`include "../lib/Interfaces.svh"
`include "../lib/Channel.svh"
`include "../lib/ChannelUtil.svh"

//module that converts packets to core data

//////////////////////////////////////////////////////////////
// Router Packet Formats
//	
// Header Packet:
//
//	    10		1
//  [ Route | Tail ]
//
//	Header packets will always be zero by the time we get them, so we can ignore them
//
// Data Packet:
//
//	   10	   1
//  [ Data | Tail ]
//
//////////////////////////////////////////////////////////////
// Core Input Format:
//
// [route | code | payload ]
//	  5      7        20
//
//////////////////////////////////////////////////////////////


module BZ_deserializer #(parameter NPCcode = 7, parameter NPCdata = 20, parameter NPCroute = 5)(
	Channel PC_out_channel, //goes to the Core
	input isempty, //isempty signal for the fifo feeding us packets
	input [10:0] data_in, //data from the fifo
	output reg rdreq, //read request for fifo
	input clk, reset);

	wire tail_bit = data_in[10]; //get tail bit

	//FSM States: i'll write this up once i fix it
	reg [2:0] state = 3'b0;
	reg [2:0] next_state = 3'b0;
	always_comb
		case(state)
			3'd0, 3'd1, 3'd2: next_state = isempty ? state : (state + 3'd1);
			3'd3: next_state = tail_bit ? 3'd4 : 3'd5;
			3'd4: next_state = PC_out_channel.a ? 3'd0 : state;
			3'd5: next_state = PC_out_channel.a ? 3'd1 : state;
			3'd6: next_state = isempty ? state : 3'd0;
			default: next_state = 3'd4; //default to idling for header
		endcase

	always @(posedge clk or posedge reset) begin
		if (reset==1) begin
			state <= 3'd0; //reset to idling for header
		end
		else begin
			state <= next_state; //ff the state
		end
	end

	reg [NPCroute + NPCdata + NPCcode - 1:0] to_transmit;
	assign PC_out_channel.d = to_transmit;

	always @(posedge clk) begin //do these synchronously to avoid issues
		case(state)
			3'd0: begin
				if (!isempty) begin
					to_transmit[NPCroute + 26:27] <= data_in[NPCroute-1:0];
				end
				else begin
					to_transmit[31:0] <= to_transmit[31:0];
				end
			end

			3'd1: begin
				if (!isempty) begin
					to_transmit[26:20] <= data_in[6:0];
				end
				else begin
					to_transmit[31:0] <= to_transmit[31:0];
				end
			end

			3'd2: begin
				if (!isempty) begin
					to_transmit[19:10] <= data_in[9:0];
				end
				else begin
					to_transmit[31:0] <= to_transmit[31:0];
				end
			end

			3'd3: begin
				if (!isempty) begin
					to_transmit[9:0] <= data_in[9:0];
				end
				else begin
					to_transmit[31:0] <= to_transmit[31:0];
				end
			end

			default: begin
				to_transmit[31:0] <= to_transmit[31:0];
			end
		endcase
	end


	always_comb
		case(state)
			3'd0: begin
				rdreq = 1; 
				PC_out_channel.v = 0;
			end//just ignore the header data

			3'd1: begin
				rdreq = 1;
				PC_out_channel.v = 0;
			end

			3'd2: begin
				rdreq = 0; //don't overfill fifo; hacky fix to delay
				PC_out_channel.v = 0;
			end

			3'd3: begin
				rdreq = 0; //don't overfill fifo; hacky fix to delay
				PC_out_channel.v = 0;
				
			end

			3'd4, 3'd5: begin
				rdreq = PC_out_channel.a; //want to start reading once we've been acked 
				PC_out_channel.v = 1; //pull valid high once we have a full word
			end

			3'd6: begin
				rdreq = 1;
				PC_out_channel.v = 0;
			end
			
			default: begin
				rdreq = 1;
				PC_out_channel.v = 0;
			end

		endcase
	
endmodule // BZ_deserializer