`ifndef DESERIALIZER_SVH
`define DESERIALIZER_SVH

`include "Channel.svh"

module Deserializer #(parameter Nin = 1, parameter Nout = 2) (
  Channel in, // Nin wide
  Channel out, // Nout wide
  input clk, reset);

`endif

