`include "Channel.svh"

module OKCoreTestHarness (
	input  wire [4:0]   okUH,
	output wire [2:0]   okHU,
	inout  wire [31:0]  okUHU,
	inout  wire         okAA,
  output wire [3:0] led,
  input user_reset);

parameter NPCinout = 32;
parameter NPCcode = 8;
parameter logic [NPCcode-1:0] NOPcode = 64; // upstream nop code
parameter PCtoBDcode = {NPCcode{1'b1}}; // downstream traffic with this code goes to the BDInput
parameter BDtoPCcode = {NPCcode{1'b1}}; // upstream traffic with this code came from BD

// soft reset, generated by okWireIn, or'd with user_reset from pin U10

Channel #(NPCinout) PC_downstream();
Channel #(NPCinout) PC_upstream();

// sanity check
//assign PC_upstream.v = PC_downstream.v;
//assign PC_upstream.d = PC_downstream.d;
//assign PC_downstream.a = PC_upstream.a;

wire okClk; // from okHost
OKIfc #(NPCcode, NOPcode) ok_ifc(okUH, okHU, okUHU, okAA, okClk, PC_downstream, PC_upstream);
//CoreTestHarness #(NPCcode, PCtoBDcode, BDtoPCcode) core_harness(PC_downstream, PC_upstream, okClk, user_reset);

// leds
//assign led[0] = ~user_reset;
//assign led[3:1] = 0;

endmodule
