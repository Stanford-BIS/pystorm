��/  �IUDZ[�d�ޔ���r��,�:vt��S��lo�?	\���j�Y�B��bF�Ơ�K���X<K�X��.��[��B h��=�?0 �P��R�n���.&�(<�L��3��r�	�W���ي��T���W�]���:�ok���JSy@�����-:_ i���]����ǡQ�K���~W���v�Q��5�SJ����,����k���o�6Syygs�eg�g?]9�	X�!�|���#�?����]EvS�Jť�K�����}	� ����P�z�nF��:��s��PN�Y�x�4�IY�yF�&9��T����,a�M���CŊz�i<�T��`��NT����li�d
Q�ĞL>�'��n�����~���"��q�l���GE3of3`�rJ���Ӈ�^�K@.ȮI��Ԧ ^�^����>���9�*��00u��qK<ٟ��g[���� ���]�o�Z���r!<�3���7�y;�cV�:z#0X�-ӄ���\6�F��Q�Y9K�n��@��ԯh�!���D����c�!ƿ.݉X��I�Gp�B&z�O��@��S!�f �;.J�\Q��Qǳ�T!�P��ؤ�_�W�!��J}o��5�������`�����39���5�A�9�s�H�W7�Fu�Mx����%{=4-'��F5V)�؛a]e�|
/!��c�$q��FR^�8��?�Q ��ѷ`�"Ȗk�'�U�_I�K�l��UuF��#�����zk�1W�]�~{����"��*��Q
Ԩ��33� Ηv��.��������hyٽ�����IOQ%�[�/{������ٯ�{�o�ۯz�L����!��I!�b��,�b��?�<Tp~��ʹ�@��
�E�Z!D�y �-^�m"�gܦ��сHz����
cZ݃��A���h&c��:���G1O��á�~�ȆNo���y�Fxq@p��h�����
?�o�oCv����9�Ɲ�d�O#Q�Œ"����n8��c��iV,�[m[F�pg�nK?>�Zr�/�ø�u���Β����H���QT~V),�� ��w2��� g���d��/>%�����"Ac|:�U5@Y�E��}���9e�`C�Nb���(/֑`@���]�!���yM�.�`�?K^q�sj�pL�7�6l����9�z&���[�9݄27���;y�F
x��T��0�~�5��g2�?�����;��0��%�\����VL�گI�$J^�`���T�?<@��ꅮ~F�9GÞ<��Y�њ��>A��83�(��
0nൿ�Ge���m-y�o@�bG��1���&���( כ���r�����"���h٬n(�ٵRe�3_w��ěo³��H�$'���;$~�Q�Pb\�����c@d1�����Ȟ�Ƒ�:nB�h�*�M��Ȳ�޲c������V��ba�E�5�C�(|곍�K-C"���Bx�e"�mk���4��}S}�M}�IuX�������Vk`������1����5R��so����Hr��m�6���6b*�y���t��Ic7.mU���W�V�3�� �"`�AGW2�(V�/$sQr����.���^�9�S>^VAK�%G�OI�)�����GN��0/��%����`Jl>��N�ؿ{َ��f޶����3�{�ԉ��_�쥕�.��Ʃ�Pn��ޝ�k;�;Ω�8v� I�6~���y�r�L6,z"]*�`������Jo���٭=5|<>���od��F �>О�?�d�aw�6��z�C�v�W��4��J��!A9�Z�5�'.~���e�c�&�M@G�*�����G��^"��8�9�7�Jd6M�4N�+����$�lG	+�K�5Kn��C�K�VzFE�c��xݚ����&�,��[Q��7����+I)��@y%q�&�!hZ��s���e-Г�w}gv��0�ÜH>�
L|�-b��~-v��CF����P���e��$���d�v��͞�Yȋ+Z^h�#��7H9.-�-�,��P�F��{�
~��'�����NҺ)��yuf.+l7��u��{����_{""~!T���*�f^A3N-��k3+�|T�w�x��c�8v����u���rI�	��!����/V����֨�\B�E,�����l_�IG��gr�/��<Ϩ'�Vr��.2��Gf8t���'1�J۵�E냅䧥�� �)�Qر}���Hs�s��l*��~�fR�����~A�S�um�*k�P�df-�>@�T��ĐEE�$���b��<?[��5vH���MH��c��R���6�ⵊz�Cdg�CW��g����e��l�v�F�G��z��V�WH^]|@.�t)�+,����4Ex���irW�'����)( R>��:�e~�a���+�+��K��X���@=��r�TR���Z�A{M�}�����P�r?�� 37��J!;�Gr�G^(���T��4�A��˻JԢ�kcc���t	�_1�ȑ�.g�:���-�}}q�{�O����|�� 4�^�a'�j���N��p��:�h�� 80�2ي���5R3��ؙ����v@J� ��a��aӡ Z|JKߏb���� ��؀��-я᯴��S /Ő��3<��x�Գ[,Op!����4c$����5`1/�����S.���d�����fd��X}�м�:�m~7l��y�oy�d�"t�Y��
`L뚁����������+ ��̈��,�?������#N�%a �X�)~o��Ka�L�ث���>l>*fc>�F ��
����pG���?q�M�εN���6,o�!������'�)����+�`�U�b�U� �C��L;+�Z���b�blǤL%��M�"�^�HO�_B�`L=Cŵ���\w���}0����ǩ ���x0�yޤl�'5�}�	�#/N�<�v;�b�����[��mˋ��傩����ɂ�FC�_~���&��^����+���u��dH���y�ˇ+i�	���iՈ���2I>>�%�nkJ��S4��˿�;id��
	�y�D���:��V�!5��0��-��J�eh��b�dvA��\X��,�I�'d���I�;^Gvrŵ�g³\-���a[־˨�՝��@lgM�쬹\�̬JGqY�������e���˶�$���������-Z�s���"<�9����J�����Щ��GQF���qv��Dh$���i�nMWcU�r���}��°�狔�{֜���(z�#�f���K;���i�:k�c:%��|3� �������V��W؏��MnV�{��/�"+����%K����xlS�D�o��Ŕ�L
2�}�%pͩ��PL�sa�ux���� <�]ׇ�<���?2<zrY�:����:p�'J�	�R�7߬l���i��vL��x5~��R��/�C������0�z.�3	=}�^Y��-Ώ�VW�E)��n�(�����-	�	��rlW�HQ�%[�!����FY�P�T��샽c��ĕ�v����� -��\J���be��
�3mt�R��(p�����y��z˸FI��n��R�\�Jw>?'���Cm7i7���[����w��B����c�i{F*�]��C%����6�?w�ר:�Ǳ��o�.BЕ�ʇ�\d��UUI�ʀ���^�
��o���b����pl�y����9�T�q(��БfP��H�ŕ���]WG5���Dg�@�.�e	��t	�`��̩��qp�y��9��|���Z7[���q����p:�pg�Ea�ұu�R��G��:D6@���΅"��wS��W��X��	3�]�w�z���6QQ��VdIY��l'fv� �q��A{��=|�B!�" g'�� θ��.r�e��%�/�so%�A�n��sJ^��K"�����(���љ7����^��=���%�@'�6T�̐���܎ Ҷ�$d8�R�s���qٰ�Q
"'��wzZNFD�,7ڑoǂ̏f���`k�j�?�����G{����uv�lS^W������U���f�]���_PQ�����]��R����)t��,�8:��(�Oz��s:�陭�bJ�yf�jU����sH���573��f%��pn]~��@��5o�s/��w���������JZ�����&�87�}1���&%��,���&��ԏ�C��A'�jY�hn	1C<��X��&+Aұ����o�K�e����]T,3����e\�>�İ6.���O���7�y��G$�����K�)�<��8������s�*A��\_�G�*/���;KF�u3�Nο���@�c����8�?u�=G8���|�X����*�����K�o�è�G��X�7b=��<�-UO6V>\�z�K�=�)d�&��<���X¿���E�bd�&-����L桧�9aJG��5��%J�cU\�	�}�<T��bwz�U_̪�;FͺC}��K^�gV��xp(gt���ܣ��-�#��.��1��.���|�ا���K�M]"Sg�a�=�͈h���uz�p�7×���'`�����f�S'�|� ��[�3�lA���N�~~YX�m��ֺ��3e�;�W��|*#�n��)�qbN�*J�]p�$]�&��Hl~�E���K�#��&f�{yJj�w2�n$��,j�k� oݡ���]O���T��\]��sg�S+�)�q���Iw��G��̐
w���R�z����ď˪io����� �n��5H�j)~�r��eⶣe}�yFa�V�p'd���E�3�ֻVz+\�TT7�٢����M'LF��"
��{ȗHn5�@	-%����������F���!�nE/�IA�歱W�@�ů)�#��)��%�~�"p�P�ݠ!��(����J�u��-��W�R�حY�y��� nn.6�<��֣C�<�Zڔ{�0���y��GTv9� �m�@��lR�ӘF!�&�c���ژ�v�ҫpc�k+~�(���b���H�B*	(pN�g�?�Ծ#G��f�C��ϣ���f���
$��h����)��:�(���'��[��e-��)����$�D�%se�|�2��
�ώd��jI�4DN5��D<�<D�g�~���B��B���Y�8��ߜ(�L���!�=��u��H��$7�.a�J�n�6�P-fI����	�2Ix�g�/�������c�,
�87�o6db�t���1���i88��?�3xe5@�m!�;Ȭ}���<�#eu)����J[�J}���K[)%�{ie��xݥS���V�l�Fz�fs�~�ۊs�H�G�}t0��U��֧��/�In.�1{��%ҭ*B	��R%2Q��<�������G	��C"�NVu8'x
]2��0�$J�'E+������- �ǉ#�uFZ5����1�e���2z�~8���BT���4r��a��H-t�����Q��@"$�'�X]��$&���x�ٔy�7@e�P�l��$�L%4))K������~ܤ��4�D7d	䵞&RG|E�����kwG�Y-¾�S��w~��'.��%�e��,ŭm�/��'�@O{�T��)�E���bd%&p��Н1c��1�{3���Q�Se��Y�z5��j���ti�������l
��V�L��/��?�o�>p�v"���3��n�9\�����\pD��d��<���Z��<��]>�yIХr���\���A^�B0��K`�'�*�`�g>RKS�:��)�n��z؃�j���]T�\�k}��_(�L=ѠΣ�X�����թ-�������	y�M�@vP��_��^=�ԓ�a$Ռy��0���m�a�������U����a���|0Um+� �R�0�{S����|k��?#�.�^��d�\K�K�W��R�~$��U��
�]HD�'�y�,��1hR�!e���;����	���Ā͜{�$e��EP�&z��֣�~���SȚ��t�e�,�t`X�z?=
�P��z��pV褅�S�����;�P�O]�r��S�����@ʈx�������,��#}!�t��|���YZ6l��s�]���|��}�ls�Y$M��@4�=f�<��oQ^�Ti
��L�dWC6���9оMs�����Ê�?Q�1y��Yh�A2<�>j�`�W`�wX�7�J�3#�� ��� L�oI��29r�}p�h�c�̬��♛��}��~E��SF;L(%�l�9I2��M���; >(�W���ޯ��ԗUF�:ѴN6�E��L��������pn��ŭ����UJ4T�/���G�u��@�;V��8<�:�:�S@��b��]��4���*]��s4fiϔ��`�h�Z�3� ¬�u�`ל�|�2��=z�߁H�G4}	���c��e�75K���I׾�mx�暦��]���W���k���-�>~��)�c����W����ɦ<����
5z|�K{`O�^�X2x��Z�X��������/�~o����[6�7SMIm�B�-��H�7`k�_�Fֆş�jj��Kݯ���뙜^^�+eݼ�|Ї�-Ͻ�<�#��1��������첛Tm��e��"�����T�W`?�b����dV~�����H�M��W�o�4�ި��BS35�\H�t�]���`��B?&��]���v��Z��*?�A��Y<*�fn�����Ě8)�..��O�4�f��g��V�kk+�(�po;,�g����7 �2��Y�g����s��[oQk+9�dˌ�~��m��Qi�����P �F�z�8� �(ZTn��i��KR�y����|�kH�<I������ �*�0eo ��{��~��Wg���v�u����&y������X�u9�#4�ʛQ˱Goy �\�E�0Qa����g��
P�,�	��{(4%3c�P$���][%�r5>f�h�E�C�5�0ӸI4��0�I�.�s��C_��PծҸ`��oUѪM	�!�%	�����a�F���w`9`u��=L�&��W=o��>
��F�N �*�q��|=8�|��F��pb��[s����C���VRM_�pU*3��_�	g�L�i6N"���Y�,V��& B��ೂ�.�b?��6�5n�NO����G�Bݶ�Bȵ^�������P�Ca�j?�˛�U�G�΀��4�6[�9)��;����hU���~*�4�lb��z�?��sW�*������ж(�r|=�l��6q�b��1&5窼��u��������H��&8�?:��N�%�D%�����a��I��r禤@��kΦr�[u�f�u}���������p�1C�� �Ʈ#*�;4��&kOa("��w�[vZ��}�E�51�'X.F�A��U?S��%����0������"��S�}Ûy�S�Q��F �w2��{V_�eu#�5�P�ٲ�T�[�TJ>��1T'0;�Vh��7��e��1������3�N�R>��M$����VX������m���z��eN���sρ� �i��vO,�h��c;%����go�L1$�B�ۓ8�3�M��]V�g'�P��[I��� /)7E{��΋T,�.JM��j�	^̚�K�=�{�-i��&MM�0.�n7��r������Q��_�B'*���f��h�$p�b3C���~\N{;RV�V[t�"C������2�	��eț��n�A��#�U��`�"���~�w�0��3����K���Ja��ڔ�i�`-�$Ԡ�_��=��r���E~ZQ�*N��|������v�p$]�Kє^�	W��g����c�ā�e������E���vO�g���#*�S��s�a�R��a��0˹K���T�G�x�)np��6juW��2�s1�⊷�~���b���j���ݸj�b����뜵z��
����}�CRU�K�!r:벹o�![��6V�U��짝��Đ���*���5J�:п��'M\ֲ5N�.Y� �w��j���yC�����O��V=p������g��R� 9�h���<��/�A��.1ҀVy���U���sR��#�>��j���i� Jx�`�1�'���/ʇ�iHs���f�%����^��h>�T(,&L�1��:kG2h�}��?:i\��f�o�A�ȷf`����� �Q�Z{�`�Jtb �6���M��x��Go�E���Z Umv���/���]�Ny��F�JL��4���ڮ����Es]ܯ/�H^�!�i���i�j�B����l`�7�%=PR�DK����� ���(m��N1��ތ26�>���O&�SA���v������\�(C-7}�k7�����<GxW�S�������ͦ5ɈN��=��t}}��q��u�jP����\ո��&d��λ�f0��4+D�\%=>o5��5�Pt�{|��x~��V�a�n�ٍ |5�F�������<һ��"�=_]mJi/$i����I|q���"0�m�}ݏ��<\���D�uĠȯiԠ1�>e�ʹ
�7��W*@1��1��9��3�})�\6%\���T	�Z����c�v���)0�6�P����߰�}��t����V�U�E`�u�:�c��|lV�&@us�
:���7�%�AާQT��CT���)~�Q�$m�ά8r�I!�$zxǽ{���@��/����U��߾�MϜ�օ 쁙�u��X���Dh�E�t�,֛'�����Ո�U�j��
O��7�=�����W�2��S)[ �0i*� �e��i><@�p�jN�"kw�g ���r�'�WL%w�/;p^������A��C���L����p+O����-7jW�bj�Z!m8`p��H��iጂ�>�E��j|r3q
�2����|�Or"���?fi�d��������x�/��^0�r[�Tٚ{B���C�a5�e^�886�T�l�왾$�8�(�@�J��b>ݣy�����hl2qA��MI\�b�P���8Єd�j��~���b|�τ���]������n��)Ţ�1|
^�DQ�y}U���,>�t��	��iƞʇ}TB�ې��K�̿��st��]5���NMA2�p�<��y��˩��6�Q�yñ)\Ҍ���&�#�6������p�մ�i@0B$�T@�̰9����!�;Jőd'܎_*>�giV�B����sE�����̹���{������0n0��-@P�v�Ǽ|X�Fa}pX��/�v�y�e���x�c}�G�^Y���_ q-RY�0O�W��Y���W4\����6�~"]6�$]�d^54����}�Op5���Lx�@(�m����]�Q�-*2�28,�rѥj��h
��C��smSE��Z�"�׀�~�Eckξ���#6�3M�����쥿�o�r��ʭޘW��.�w�9��^��4���؄�������N��o����g5�����E�VgE���lۀ~��*>�7b��鵧����{tly�F9c��z�=ѽ��߻���-�mw_hy���ܶ��)D�-�÷9�ibn�b�#Ċ�B%�_1�����H���A{�&~YW�e����%B���߃@���C9�&�`S�������z�i��M�c8JN^78�"��ŧ[�R���G}Hy�+1/�
룪a��ٹ{����N��>H�2���7�y���Z���<��p��7���x|A���w�1��;e����4k|�]� M�f����������x�K�&|�&X�N���)��S��t�aV�7.���B8'�>ޓ�p�{��X�θ���b���Y��Ц-��Z��h,����,;���8��NQtr���(G;վF�:�� �=�_<AX�|O�
�I$��~�٭&i>p�=.�t�]P+���~*�ڐ$�0tm�,3Ϝ�%��Jw���GTB%�E���4燣�A�W%��"b&�@S�(i����H�2��BW��9��<sa��۲�1/��Wz��b]�lH�����f��C.X��o)��l.N�j�C���kyΕ��D���ѱX��
�S�~#%���S'�+hXj,A[�63�cu�0.X�����Q�U;�(�y���30��-5,|�h�����C��8hb1��RH+j.��80߮�r��n����]Q->��52��P�PVH�b��[^���z�i��̈~	@U%�%�{ܛ�b~Yh�B]&I����\T�}��R�g4̅�K/L�1Q��ASV(<)m�~kQ�w�g1�����M�oS��� 8�ȓ�|���,��.W$�l�y�vH�W4���g�&w{8�O�4�k�"�}4�yw��gd!<6�1��G��|���}��r��J]c��H�M�9e�&����ɼ��y��������\�F���N�]��/��5�`n>���������kY.M����ܽ��-B��ES��E#�n@Dg��M�ܔ*�&�/9�U2�@d��H������%X�>��1n�b��LXC� �E,��KSI*J�ڻ|��眉N�%�X�u0�+�%��M���3og���8�;H�>��i���ֵU?LM��<��7���Ů�T/6�X��Cb�W�Dwĕbh�t���8��y�(��)!�$��	���Ɏj�K#F���
����L�#�y��%	/%3N�1��g�"-ǽ�Kk��+���)0���@��]޷�E�ެ�|k�I�����:Ec�$A������D�k��ţ�.�IF�I�.�(�(5?�<�c�3z�ʢ}���f��.�3���Q�"lm����`�0���S֔b k�A6�Y�אg�>�kO8�kg��B?V?��Q�{8_��!Yr槐��8j�ݩ)�!b!Ӧ�\����u^a��,�ٻ��2~�r�(���e�=�^��T� ���%doȪWqA{F��?k*���*��My��-<�R��k�)�������w�7�J�k?�UP`�8@e��8��S ~ך��Q&6�R"�����P�������>�p���\��9��R~��x-x\�\ߡ��#y��7@��
�ۉ(!!�2d�f�Xyi�*�3.:8�����1�If��P޸��1Ehyp��fe;h?���$�GOfҸ"�c��݌��e���IƷ��ڷe�ϷB��\���i���T�'��\v��tJ�(�Zx�|	�˽��fMr	/�T��&ђ�N� ����G"$�k�h�L��|9����à#����_8��	��=#��VƳ�kՔf�Rnp�oF<�OAN�$n����:�Ô8D��ȱ+�#��Ӎ���+�����{�GY6^�mq*�n@[�1}}���F�gw
�"βn�]���΁�r��s`)#�B�z0y�y��m����U�nK�5�>� �$��2�� ?=q�h"�"��1�p��9^�~�����ҽ�	��y�2�JtqF�D����`�C����HQM��>%ߚ�O����i��d��w��-q�F�	"�� Z��lc3�F�Xi�+��,�ꃪ��������w>W_��mQ`�U��˙3�j�(�����ivؿ�Z�J+��
�l����F�0���)UĄk��^d�Jg[V6Ci��4��Yl����eP3�G�H�E>��F�)B�YƄfys�/;OaP�A�|�~���9E�/[���]i+^��#]s��{�N�����Ƈ�L{�s��y}<���2P`�dS$�L�M�ډ岽�-A�S�#�myT�gsp��6�)P{Hl�1�Q7��y�!�X>�?�)��ŋ6`��X:�σ�{��L׶Xo��V�_�^|S0��V8����P�e���R٣� ��O��0� Q���ں�����9��߮��|BZm	��:���+�Ro/ȕ0�G�]7F�x۪+MS�Ǟu��$�hƴ��e��W��@����&��!��D>}�����q�p�.ű�(�C�����hRBjO�+���♄TMm0.��J6^����iE�bQ�gca/Bl�+D�}%ӛa�=�h�Hu�����:��b�-��.�H�(�TY�����KؔM�B�RK��0�sѳ��s�[��{�Dpy���a������Og�h�dK�a��vt����R������[����,O��a_{<�m)D�"[��k���9a�E^32�{S�4��Q~���+<"��$s��Lݶ��1�fRу�&Mض�W#�葳�V�=a߰~w&��=���iOf�PW�=�����kw����B�i��12�T�eE8�)�0>�ttH�=��_�η$~G�ʥ�H��i؅�6�v������ζ���/�ۧ�
�&���|�$��ᶠ7j���I%"!�l��̹��)�P�\�J���z�GF��P���y��;������k	�4aO". ��ٸf����C"Z:�6�{���<{ϣ{�	�'�4����*wc5��y�jP�A�M\�N�fѺ�ϡM~EG�Nw�	 �R��-��8ʱ>%���t`�՝�x���!kCh��b�-�.)��oec�����7e���6Q���̟���|�m�J/-w��8+F���v
0t���0�u�>��s�r`c ���^�"������>�'\@�]������h ��NY^E�$X.��#��Q]����F: �:{ 鯔�&���D��C�\�ߑm��������#����*:J���ɼ;�Q�5֟��_|�`��D����<�������W����!.�����*#�i����'5�Z��r�R��eg���nh:���\�hq��/|��2'��3�4��S��N�򻚼����7f�px���_r�TD��������kILb@\V8}m���X�X5(�]���z��p�
�<LU��5�Gˍ��g��M�7ɤ�Y�2:�=cM����=H��$'oy	�ȳݛ��s��6�dQ�J���e��`�b�(��@�̱���7������n�ܝ˓�:��&��ϪNe
y؊&����A*���ˡ�aއY�9��5�+;�e�N�?�%b�O�d0�#+F�n��or�mUPg�U��Ic����3\�+ �a��R�jm�����T
�;����}�0k��Qq����0N:����ܿ�eu�8g��� ��ǋ�Z`<����f�V�<]Ȉrbɾ�0 pu?�<WT�i(A{u��2C^��i��ho�yguœa��'A����,�J�25�MюT`����<-W�G{D ��!P<�p����Q��D���o ���Yh��:�(%u�� ���,?B|8�ώ`��m�s1��h ��'��΁��A�w��o��T�<df���&��Tދ�B��Ԃ|�6Լ7�YǞ���Q���F6���0YRo����-�+�^�t랁jk��"�ț�����*}�Rʘ=�8��P�g�m��ҕ����ek *]�%�8��k�ET�tq�!��rq`D:���Ʈd�ͷ�"���{�8!`�:�����k��
h��p��5�:���]��+\�r��4��#�%O�w;qE>8N5.�ڝڨ��;)��o�*w��dn��t\�#ߦd�����^z.&0�XO"n��26o}n�0 �������,�΁�~��t���\����]�ѻ��'�H���6��Yb����i�cނ�Ps3�}��*$�ܴ4�l%P2�t�c��S=��yiB�ؒ�)]b��Zg�'�� "�y�~A�(P)z�E�l�}l���!m��G+U�OR���� �| v�"̢�14��k2���������e�X3��m"ӱ��	=A->�Ĕ��z���֜Yd"�8�Ԯ��?s2�
�u'ɻw���<�AN���?�Fu��ۻ-�8 �.r2��	r�d�G�
oZ9w��Yb1�[lp�����v�ss-y�^y�۵I-"��x#{�1l�Bg�~�l�=ɭ��sՆf
�fOU+��X(�T[1<ڰ�����?z�-qUebt�2v멧��7�]��g,x�)Dߗ�����R�N�ǅ�[>#vZ�:�����N���
�bR��0cl'���A�3V�<���>\:���0$�i�"2
5����s LUbΚ��[�ޙ"�k�0E���K��;J�.�Z���H|̒
a8�DX����?']S�E���e^j������%��C Fk�Q����$�%f͔�#���u.��ݠΈ3LWiCf4�����eV8�������`N������	���eNib�#���oo��ݣ��3�}����J�W1�������&����Y�s)]�!�9��7!�n�OXI�d*8㫖t=}�U"�򾾱���[w8$��}�bN@����<�6��ۺ����
�n� ���F���{fݎ�(
@�A��<)��j}S5h�Tܠ��]Ұ��rʌ�.SԜB����e?e{�聇���~���6�z�ֻ��ܨ��g3>��ػRٵ�\�4��L8�Zj���a�T�o5[���47�[D=[�D6X�ڸI���?͖X�Z��}�"���䙧< !�O�P�(tiA�x�Y�9Ѹåf�#O�sɖIP�r��C���w@�^�.�����<a�n2@�/��8�Ŝ Z/��8I�<{A�.?�~Rl4�eJ	X�w?J�̫9Il^k�, �s�P˜^X��u�O-�u$>���:>��A�I��y&�x�0C�P1 �ǔ��|J�r^)M��y�{K)���\ʋ6<D��!�|ɵ�+���� ���܇�a$O
�M�Q�������u���_�`Te#��e((#5�8BMl�DK�О�����<&�O�+���8V�j�7]�� �����Z�1�O�W-���tF}�ՙ�%Z�;�ʜ�I�T�c�\�ZwGr��������o���C�BQ��:\B�C�3�+�uZ����H<Od����Ϗ��>��1��w�]���b����*񃁥���Xk���Et���������t���*R��e�Y�������4`�˧R&�_Ș�)N#�L��W�6�����u�iY�sb�p!(ߒ�^�0�{�>^i��+�gv���}�z�-���_t���|c�|��
�����O�%��=Su$�l�%�Q[ą��A����!��τVC����T��֣�7Dl��'�hx�8�>��60 �N�GY�SЩqjx�PY@�t�%{\���y#L�n̗��$6�|��
�ųc�I����#�2<yLa�ol⡪�wVp��M����MMI.��ݛM��p���z�@���娪�0FB�m5"��RD��׼� t��1P�Rv���K%�5�����Xi�V�Yirk0D�=���������:�}�o2��$8)T1�2�C�M��?l��0��ٲ[5I!P�DIR�a�i�ο���|� *(��. K�ߑᰘ�Ȥ��1��X��#Ì�Ye'��ъ��������\����n[I�D�M,���Syx2�����,8�CibJ��D���� ����Y�a4��Ө�FU�3	t��O�W�Fj?�v���J�dt<�$P"������S��~r��1.|�u5�f������.��@b&����~��D�����O��U��-��͹}E,�V�i�Ǎ�'w�<q�a�jt��4q:"n���we��J�34ww�z�n�I�i�1'>���u>Q&��{���p����Nn��L��hD�e@�$)��l�6D��������v!t�ze�n�xu'�h��:�������+�{$]�庬k�5+ X�#�יܕ�jS��������/B��b	/|m�8 Q����쭯���$w�������j7(�Ns��:���(:�M	Ƈ;�FaT}�?��7��jEeA�g?Y3Y�^�_r/86Zp���S��c� 0S�Z�Dg��qxI��X�ԉO���)�%�%��=�� �ַ�����4b�+�����V�O�($ߗA]�<�V*���Z�m{��2�tۨj�5'��Мu =CP�%���T�(��Dُ���x��\}\�oپ�
���M64Q�郄I؃�D��9Ca'��:�#iO/<k���!Cp�~�)�r������a�+�����_�_�T[uhN]�r
jp6�?y��OU�#c<��;<o�X>�ÔȺf7�B��a����+���O�w�&��b��H�S8��E�-m{A�����p�Sn`�:wPY�b�����W�M7��F.#�kp^˹���y?���⨏�z�4�LQuնb�����=@P�J����5��;�C�zZ��0�>�lv�rl�Pу3�����m�s�X�� Y�Q�A!F3�}I��y��݁�3��H�/@qR���#�Gs�
�!�����\��˓�\s$��;
��G�*{i�_YZ�ͱ��HR�y�����k7ɼ�m�P�e��*�:fF�B��kaaQ������@/��V~���O	PI�e��Z߳)�y"zb.&�h���+�_0�5F@m��"4�g���Xu����ww�in��y'�Epak5��t (�Fp��䛄jٙ�&��6'�-C�����Ě�hay]�$i�9�	QlD�P-�w$֌�>�z��J�\q9�H���*�����J�)�dEC�c��Y$)u59ʸ22>Պ�f�����E�W�cU��X<���K�i%��G�/�BVmq���V	5����p���u�����'��`>�SB}���p��]	�I��Y
Mzfl'�i
�+k���M�qN芚Ek�w/S���eg� oP��[ �ye/>D0�����Q�zɃ�6�����v�r6��s��i��
^[��ۗ�q1RJ���I=Of[at�)��?��[��;~�so��3�'�cڦJ�n�|�;�c:Ҕ6na	�:�z#U��H���<�7�s�{�wd��rM�_"�#�y���4�0'On�!7K����K:C��i��Շ�ԼX߼�����?(�%�	��)Ȋ���9����N<��flќ�fzA�D(�&����2�N_BD^��N���\�����6/{4K]ç���y�L0�����3�o
��(.�.�~${J!�J��x��5"���t� i��X�&	��S-�Yx/��}�h��8�:@Um�pb��|��z7Z�+Z����R�|pP@<�l���=��< 
�]����]��������'����>�_g��� � ���K�����QR"~�=f?|>~���:���=|(6��N{#����VGM�y�gw:�*1��	2�V��%���S�9��a�W����C`t����L��^�&# �#�ʩ;J�J�Ұ�LP <<�5�e�a ��T#�h@a��	�9|�������/��u�"bA��X�N�ïc�kեؐ9�ߡ^��ѿH8z�i�p��p�4��(�*�T�/�=eUt�[��r��'�������җz��  oe!��a5�a����l9t*'V'��~���tg�pk�k������9�M�ֱyO �JEnEv�g�fBiNz]��H��	`~.��7�(�X�[ۢ��w0Z��+1���_.�\���p�F>Fs,D1;��,�xf�_qD��T�R+�x��OVm��j���`�U��7�6K�~m5T~z���D�Y�V�B\��uH�O6�Fھ��y����C�؎3�`cĽ-n����5���A'�q�B��~��<���}/���j+�P*�n�R�&LP!��}���O�r6�[�C ؿ������\�j���	��PcEݍ�*|h��]1�,�䥪�B��n��6���歒�f�F�XG�؁���[��PՊ ]IH�׾��%n�P���rj�pg�>7��wi�{�ҽ�+n^ﴮb񱤈�ʔ�V���e��S�#��Bao#�Zϗ�q��Tx'֣P���↵��7�J�q�U���"�i���c]���>�2���P�}���;�J�zGA���n�?�����RFtj��� �2���d��ٺQ-�-���v�J'��)/�K{s[�*�"��x����o��������FN8�
���۶�;��.�� ��1R�ԍgƃj_&`�)kv�����	{�l.��؄p��P�W��_L㾮����#	�'G�{yi�✆A^�pC҆,v/�0(�v��R:��<$FJ�G��]����6���#�v�]f�����!�F���!��aX�浖��~�Rt����M�*v�'$�W<j��8t�-�eg��Q� �GK3szKTϺ�0������a;����{R"[�s��J0�h_�pT�|}y1.ɴ~�x�l�X�� uIk��,��Q�O)L����O��JT����ȭ��
>6�R`x;5S�E#k���<pyG��䉫bf��Ҏ����xD�g���#b�=��|�Zg��ʌ>Ӛ�"�_�WĨ>�� ��;]�����n�Ր�K�r'ɿf�v��[�hn�Y�'� �5�l<F}Я����*�� ��b�I�z��D��5���XH-W	�K�\�m�@T���)�g��z
�|K_�6�p�Y�O���}m�rm�7^]�Ŀ2��c�)B��H}-T��A�� ���T<1t�s*msG�Jv#�elJx�{��᪣Þc��J�8�*0�r���i�	�=$�#���׎7�ￌ���/�����e��JR)��j ��� ����������������n�Hۗz�%��P7Ý��U�]>c5o4���qg��'�d���)�2 �8�گW{w�:�џ�������,�x���m���B�4�J���3,3d�-'&���xA�����e��RJ�-����\����T��Z6#9������o�>�ğ�צ�A���n��
)���N��q��q�8�]Z�f-����<�D̷��h�?w�%�L�n�2En��̓���HsYc?���7�kqJ&N��H����ˢOб�N�);<`��m�����{�8b6��C�	p�x2y�T��|�@�r���b�]\G6��依��\ꯨh�@���8{I��Z�/慵#��.�����.b���1L�0��;�����%B+�����kЬ*K�Bm��b�,��$�^�Ϧ+��~�4;�b4F�d�b���w�N��2Kw�~Ue��0]Kl̫N޺�>.��p������K���~5�����b=�=C�d�n�X�&��`���;BQ�m�����5��3B���1R���2�vZ\T<Um����-Z�]ḏ��C������f��؃f�K���K���wZ�P��b���ʟ�(��M3ݼ��;F���C�����q��:���hLM��$<;�~�l|���ѕw��T�V�	E�.l}!����׹���ճeLm�˚!��b� �>�qx��%�'Ɠ�ޘf�k���s��o#1�	MR��dy�:�����!Fd���JȚ��nН��a�j�s\.c�:�}q,���O"̙*�.��.{��;���l�YUI���$����G����#�9��#i�3�������뮭z���ǭ�0�dgxZx=���d�eU����1.�fZ��n���j���\�M�L�dZ%ɧ*�sB�[v�t������u�2��b�\���v�R��-��4�k7���?�G�$EwA����W/�b��P�e20+"vD�{���1\���ɌA�Q0zWS	�9���z��72~�c�|�x�d� 09�E�ï�ِ�C7k�I��#O�/� ]���]�1���R���o��[B�:���U�&�M�kag��N?iz�Z-��|�m���-E�#}�ULW���v I�&5���'���rO!a�GD�A�(���i��6��K� �����O���a��r'�'�����&��"�ceľ��.GT�(=Z�2M�?��*��NΨ��f�`F��%�Lr�����*�ߛ�S��3����t9�;3���Y/��D�������M����!�KDo�^�Y�{|�t��H0�Xw[K�&kTy~�6H:VG����xd!cT-�%�~6�@����AӠ;k?<L�Q�E��q!��/��6���..��7��"9:n".����-�!�|C� %��xH&K�wb�.
�VE�榧F�p�_�4�3���L\���f�s�k�&c(�r��%y�i(�����ٓ��оId�(ҟO[ӷ������2�m��Γ:�Q�-�)8��qώc"U�}ۇd��θ�)|\"
�bQU�ب��i)o��@{g�n	��l���5�܆��!�`4词"��	�����;��(@����`��d���yP7�4z�)��[A�
�� �<?q�b��ft�xZ��ƺ΀��?jV���Rp�M���2f{F�-�n.�k>\��6���`$z0���k���*�V��l��������O0�<���h-h��'դ�+
aPJ�R���ڽ}��eW� g�:CNب��!�+Fq��&�@�no� �W!o[.�X`10}�2��?y$�(W�ͩ�.�\�z9(�H>��n�m3����n��z���a�JܟO~�;l��.#BIJBw�2ߖ����/O@�"�r��d��оCs!l�܎�~��� ��-�>�7uG��Y���đ�[VJ����*�'�������|�W�&�Òv�*�����'tu�o���*]�ރ�฽m��I3n��[9�c��g!0|ģe�;/�l���ӱ>�|f{���ߝ�cvR�I���G�P�I�"���N�L=��CH�n$ı���A���J꜑f�h'/ɴX�� -U�Ӂ��|�\<����(q�fv�ǥ�����E9o阮�$�)g��=^��y݅�v�)������\|�K�f����p�6U�d�%5���`��(6�Q�%_Sa0M�ŗ���4P����zI���P T����ő�a��!�c:�J�lڽ�I��n�/.�&����	e&�^/���<�O�����+����I��Nf}�����F'��5km4���wm[5��Y/WIMbq��2�ޅ�8I%t���e�z���9��06\�=�� X#L���r��S�T��^�$��~i(�K0b�,B@��d#������>�V�aD�x]�yn�Eq!�^YC�g�[����x�*⨷��]�^��mĘ��0e�y��1{�!��h#u������ǴEQ�ǲ�IX�Y�Qn�-�^��dvT�m�`�kv�!��Y����qʛ�$qe�.�l����ɖ�������n��#�[���ҽ��h�S�� ���v�o��tYW��.U�lV�ogQͺ��1`|]Y�ڃ��8�62h͐��A/D^-3�ռ�Q$�(���y�#1����Z�U!�5P�t6����8`�2�H�R�ǅ�I;��PUE;��[wO�j�P_�J���p
�S��3��3�u����T��3��M:�Sj�oq�e*r��)�#�Qe���d�Z���+�F?Y!(9+���gH+�|������g<�p��=)�" �[$-��Zr�@~7!@xLG�M�4��*jǒ{����]�\Hz/Z�'LM�W-¨�aĠ��t)L"]�y�mᎡ��q�2"�g�4�!8�S��~K0��F%���Yާ4Tr����7��X�Q\Kg0�C��95�akcV/���O
�t�V��Ύ���Ou���;{��k�Zu�hi�j�C�|U���ڂ��˴(+�&8@'7���|�!�5a���̅�	���%d���V̢���m��������v��p�p�l�7ex+3�b`979	߇=b��?9�HK�#+��9�w&��^���'J��?��㧛܌H#�<\+�7���ت:	/�����:�63��~�ܗiK��	�W������:��S�˥���M��4�g����cH~�)�*�������Mz@e�>�f�Q�mHp^	�SSL}��@�!��Cra��A�^�m�R����.eE����CR�Y��t�1?�s�מ=�k�#Ħ�# ��`�t��g-�G��h�o�{B������U5�����E`D�8�ȶey�n�G�V�q���[�鍂Wʁ�S��d|�t�)AM�=H	a��a�����0��KZE�d����\�
\٫���C��gY��@�D�,�`�Wl]��	���><�8�Q����)���ֲU�]��0�2UG���-��֥Vʑ�u#�ҍ/��D�-DB7�����BrT苐RK�Կ=A
A3�s��m9�3�N��8_��v����Q/2ƒ���~l��ޔڟ����	d�5r IvU�jn�;����^�q)q��ކ�*.g�|SӉR�i$&�`Hgi�g�Xpő�W�#TX����"�� �|z/�~���r����3_2�F�>��P��rH~��ʶ�|z�&���o�2&�v��,�q�ļҬ{!M�A���}
�R�"�8��j�N��J�^����Lȸ��ȴ����L���CO�HD2F ��C�4�t�-g�%��dR������@�8[�ܨ��D����<̒5ʔ�?��o)�P�c��f�[�.Ȍ��+��,��ˍ���D��@�b"N@���Zӱ�*�u�j(��Ȑ���[�Z�����u5��H;�\H�w��*�2�o�-.�x���N�w@;�����A�Ŗ��;�@-ȣ, )��� ���D}�W�5����,R�0J�BJ��)�h1�F�׼�Y��/o�3�$�'���Vc�C¼�²�ܑ�@"���[�����vd^��7�vO	���Q�LqM�5pe��� ���G���^�|�&�=)�h������T�7�%��dbu���l*�� ���>�2۸e��H�^�X8 �%  n������T[���%*������A{�&v��̭U���w~��G���GHM�%��s����!~�Ln|��
�*�+d0l%ъ�������QXb@�>��pˮ��-�R�w2����e	Ǔ�z9���f��0Ѓ�O�����@[�!)�I�TRޒ隍I���W��Bp��� To����Ͽ��	��-g4݇gu���Q� �M%�[((d�n��썉ѳi3� oj�b�(c�ڼ���<`pĵҳͷ�O:	���أ�9�[;�-��j�k�y�@�
�a!Ԛ�h/��+��8v�y�D�����U2�+b'�b0j�����A����Py~Vх:xI��l��{kv��aF�J�,���K{���W_�,�H�Ǔ.��?�ظN`1O�nvl/?��h�y�Z
NAt�K�#ִ�kmf�	�Zl��0*�e'�B�b�(es r0���*��*d�Z�`��R>����@g�ued��NU�T�z�ɼ�h�����*׀�ymo��z� N2yFy0CD�jܴP�D��r���,�"�Kd H�ǔ��1m��1����r
�#M%�k-p��P�e���AB�C[��.��+:x�U��[Z���E\5�G�œ�=h�@�(ܺ������[�uEU��=	�'���4%i�qQ�!��Vǂ�q蛮�|<HQ�!�n�?��^O�k��1A#�l#Y��3ӭ�1*�ቈ���]�"	��ynF��Sm�3�*V.�Qz��13:��&����p�6e�7�~B�x7\���Zg�A��]y
��P^6$�ȃ�՘��`�k)tY�c��.���ov��M)yo&3qm�W>�E��G��,w;Q���&d��k�Olv�=�~$�{nS��E7c��b�L�)��͊X��@Ů�@p��ѧ}������6z�}9�����s��P��mBV���W��c�ud���Z�;�
��S�P�9��=
�g`�����ũ�8�3��]U+�ǘ�bki�Q�B:Gq����V|]_4���w����0�)��1Y���/�!PC�S]:��9�H?�{?��V�c�1HHD=������̵O�@�׬6O<~�����&���h����Ӏ�PBV�FvZ�E�6�e'��|���;����`��\�H?tnmY�^	ju�>A<u�S�3���*Z���a�4I�a(#?�d��=���۵n��d���/��I5�����А[��~xdAEd	��f��1pclW�v�s���b�d��L)&�	.�-F������n~n��W�nM�c.�WR��I���^碦æ��(��7���3ַ�&�:����uJs�t]�C���
�%��<��j�L5��]���V��`^������E�)#j�ڈ(�'���;�;�K������<3r
�'x����^���Wg�`/{�A�S��jl|Qn�DR>>�MA��އ��exҫt�iM�O)&�Ǿ�&[ҟ9�{�ݴγ�����]F��j_��.�X���CX�8v�fp�Q���Ď�Ie��)ͭ��2��{�N3��$���U��M�WԨϵ��g��8pR�܃�|&Z!+ʿcô���4�Ӕנ[����hEj�)�N�V�Rކr"R5z�	1��,G�&�-��HÝ�׾���t��N�T@C��ӵ��i�R]Q��v�j��a��
��f�i 4���}B����hp�Up%�.+���ky��!防�:���R�Ր�c�����#�~i��*��MR�Ҩ��TN��! y#:�C,Zt�B�Oh#�XĲH'/c�XtЉ+�٠ψATQ��r.���к3��;!�|��yPt�jktk�#��w r�&�?Ӯ��n����8��S��c2��1�?�֗W�Ơ�x����6M����x������m�#)˶a�K�	,�$²��'Tc��3Ѥ���ڌl�(���[}0�󏜮�`�!Xft*�� RF<��a�f�<�ږ�n�kl!` � ��;Qw�"?��ykQ�~P�ѷzUjde�6H��_�r12�AA-G�E��*��֫mdn�#BZ# G�jn(�/���������;md�4e�u�y(Ms��E�]���}��t�0�a�;T��	]�W��$l����e�� �޿�v��<'�@3��=.fޓ�ȵͮ��QxS�2� ���n�ͽ����h��t�"���li�d�:�O+֙�B��[GƐ@�!������)��� �����\���E�`%��9�'g�	V��}ĭE��1�� �s�3 �~v[���{�b"�*e��cߣ�|�[���9|+���גlğe
(������v����:m��LG��-.	"����9r)����2O[\8��2�f^��ɍ�uI.!�5�eAA;�h���V�NɡP�/Z�&�'��d������`fXHb�䞩�
�0�̾z���X-�0�M�2 3"��e;������x���Mt�Ǡ�?FDگ��&H)��KW,����98<i:?��v{(�w㭢���r�{ˡ�0�u�aU#	v�@��~����� i�ɨ�Nr�P.*��E��U�2TȪ����������VS�����(���^�@�I��ŎS�P+��\�-�p���x����pԴ0	��,F#�~w^H���oK�,y��]��2CI�O��D�F
���k��:U��)h�đ����n�e�8�l%�M@_3HΥ��*2��97d�9T�U�nu�n6�?�f��0�ˣ(�BA"V����o�ޕ*��4E6-2�l,L�@���	�{���C�)wQT �n�M1���K�4$���-�ά�<\�
���t��=ڬ��_���s�1A�~�{!��zp��.
��DE�����0�Yܰb�{LnᐓYs7}!c$z2��$ί�P���_�a�82�|�(�ő�2�9�6~j�.��Yi2��I�r Wokk�žx1��qi/j�2?�[���p��J��p��ˣ���#1uQoɾ���=�%Z��~������KG���L����~�Cue3���W�����_-5�Ž`/���<���W`�N6o�<jǂaMp;'FW����$��|��i�c�?��Γ��g�>GdlC�(�����'I�3�znUFs�2�,iXc�ry���bth�� b������c0��y��2b���W*]�i�I�`����>�ֵ�K&6�
4��WSx�il�Z�˓�>7O �f�(��r�\g���zp}���JQ�:��G���<9����U��Y���i�y��%7o��%rF�b����kydo�U����U���T��)����G;�kӷA��Zt� 3�4�+�ijĥ/����*�v�� �E��8Ff	�q��k^�\{�q�'<S^c��v�M�G&�4�Z����eM���BI��"����8]��r��^��*��RZ�ȵ�&9�$o:�{ �<:�@�lV1�z�I�ؗ������);8�$&h����眷��cf
L^el`�Î�p��Ȏ��폘v����u�G3�8~@%J�n��>%�^�#�.�K����?�,��Q1G�o;py���P7N��y#�Y�5�w�Y3�$g����[�ؒ�׿"TnLF"%��v�}P�	`+�^r��Eň�@1������O����Pڲ��#���h�k��Z�x1�
<՗�@���!�2O�m�Q�R3��Jh�t"��]�A�.0�j?�/Ifn[W����$�U������������>�%�1����{����S[<1����"Nk���^|�Ԡ_'�c���,R���߅DR4�nB��\�)�W�}J7����K׬����}�/T�����������9�}�K�i�43g���0�L��u�ü˫Ӗ�-�Ee�9�M�X�Ɵ��m���7�"Na+@"{N���n���*2��a��Y��dN�Ӂ[�2��1*)���9�+,�IE���s]N�t��zL����@)C1�ـ�����˺a��"Q����4'x��ɹ�g��5w��+�׬9_�I�I�<���r���?6Z��4^��
�I���<�@!ɣ|�f��:��O&ST �㤌���|R�*F��n�q*����6)�z��b^%�dC�Oa 3�)�|�}�4��[$����P��i����ztf'�pi��!s����?�?���y��1� ��wZ�k���]���X�R�>̈́0�Z�|=����	�G�j��Ǘv�|F~��~���B(�ۯ~
廈P��
j���A\8�>ݳ�x�K����T^zɶl�:�/!v�u*�$߿�1�n]��u��W! d4�6�� �'�3�@e|.A;@5�����4X4WF�m�˝$��5uI�0���$y���	'�i��R�@��J	�VOps�s�������Q ՠ�gY�H�+�A4��m�z0��Dyd-΂�y��^Mԡ6��JT^u�tڐ�����3v{�="����q���A9w��}��md������1X
2��1�GI.Vʯ8��DE�~jr����:3�n!�A��|��%s���V|��G��̷���q�����s�_o�R�Nh�`?�^#2���˄�I]1�G��W���)o�M(�!v�,&5���"%t��ɝ�^�SĢ:k�'bU��w��Op�i}oW6�#6�Q���x� [u����̍�g��p6p�&�9_jԦW����l�j�{�Sy�[��(豌y�<�+O����p��]>a���BO������<���@�lr����_�4Tu�諭��E�����#/ߛ�z�eXǂ�uUݶ��&\�2��ڮQ��Z�X��PzQSoăI=�|�LD̩�ry+Mz�dܬ���o����8C�ڲ���b���r�gњ��,��	�C�n;l%Q���{�tp����ڔxM�R����Ks3���07�b�g�M��̄��͗�k�ċ0b:zQ7�b�Q�0*6^n�<߆���h;<Q����p��]�s�;���AG�0��m�H� pg3�Wgz����@\�� ��y��R���4��y���po���
�Qd��9���-�X�M�U�ut���RN�~#o��u�B�D�+�/�or��G������[j+�h��A�t�$��ie`�̦���Utx�Q�I-*��DQ2�n��#�Ṁ[�7%�v���i�6���٩�������� tT�D,{9��=L�=rO>%������=?�i?	�s�`b)���?�!���Y��6@0{�	WZ���wJ�.Ŗ[���ډ������ŭ�i�=��ɠ�����������
z�E��8)m:\�
�QZ8���+�g�$�o��v>{V3��0	��}�^~A[��8�7�5���Ѐ��.�S=�o�`-Ǖ4�b��F�69��Ė�nѵcX ��v�Tzcqc��o�̛��\���$�(p�o���X� ����UV��&���`�x��᱕���3IB)0I���x���u����W��h�zC4�D�h�*�r���y�7����1��x�y/���T���9���X�xp�;{�����K�Q��b�`�ޯ�ᬜk;�o!%H�
���*c�g�ݖ�D�br��TM�M9F഼00�oX��朲�Iu�!���sZ�0�Π�HH�˄Y%^��A!��*�o+�7ݳnJ��dfs�TG[�޵�m�i��&�[.���y$Ȯ?> 5��D����m�m����{�� wNxטb�)+�v����
��V����*KF�x9O7��� f�������R�P6�e��6�:�O<5���,z��
����Ҍ֓�-*�f�J[bdz�8)�k_I\8=F�8�΍��M|7��Jä	'k,i�Y����$��Yc�Fr/D0���N�=1�²��5�*3+G)�4�A_2-t���A,/a�-)�2:+���7˝qmd#nDm�̥,񛉷���g����*F~�5tj�7�r\�h��H'�S�#آ)1�E��\����@� ����(���1�Լ'$��8J�5���h$�c�8�D��f����ן<��!1��.>�hEߵ*X�?bxb9ޤ!��f��\�1��}���	W��NG�x�����R�]*�b����{��ʂt�+��*����)L�5r=[�$k��ƚ���G������n'���-�i��.�ʿ�$�	�����t4�f��s,ϝ����R�aƒ=3�
��`���j<6�wՈ��os9����E҅�"�2X�!m�M��Ɯ|i~z퓞�j�4p%*�6���Ό/�}[J���x|��}�?/�w�������:�Բ@�����5r���j|aZ!�9��M����:O�g۠S��ͪ�*�"ĭ7x��z[D�9<8��l��y�'8��X�Qh��W�pF��h��i��|0�ad �5��0�Փ�r���4�$u���O��xh�T�CϏ�w������BYQx��N��~vʇZ\����/�$��.E3q�YJ��ᓗ![6s���nI��ӎ�e������eJ�M.�����}O��'��K-K-��1��%H<ћ]D9�`cNsc3�&���=����M�)8�N7�8����Y��L��ٝJ^����LG1�KzD�l3��]�iheu�r�����̘�Z�Z9a��?�=���:v�{ t}�.n�7�o�/��C�&x�&�|�Eo{��P�'��gZ"`��i�R� A�k�[��d7�V�d�����vՆlEE�N��k���^��5w�ϯ��# �e&�q��$w��O�U���<���n	2�G�-��ފ������a�=���J����%��A�x0�|
�r�W��.��+^�����ϊk3џ~��j�
Rm�4\����/��z	A�3X���k\��2BYM�A���TI5�!�g�T��c����V��Ep���K��������hq����LѶs�x�޶�)dmR�.��s�qG`*��M�%�<g�=��x�uf XG�	��K2�5�&%/��D*A�w�aa�X�|����4/�q8�4$�h3/*���޸���ye>6~mV�Dy�4�ze�A����0��qhG9�쵯�����ܽ��x"jѡ��~�j{I����(���)��2fA>�l~"a~r��j����&	���,�i�1�B-<�ʎϢ�0A�}��9{�x��R�f�c�YLL���m��H0��*�G |� �@��V�.:3P�5b"!_�LkL?�ݼ_�G?W�.�wU[�5���%�K6��d����d*l��2'H(���Ƚ
s���!�L�ch�&F��)ӥ7-�w�Y��U`�=��&�
]�sΘ��/�(����y��������j��X{�e�t0����Ӝ0؂��Gl���EykOA%��،�y��7R��b��tzpvf���7B�i�(��$w}���C�oo`Ą"�M#1Q�,z���O�7��A��q0#��!�E��q.=�+��,��+�Q!P]5�O;waÛ�`����.��7��j�o�(B+��J��n�k��)��E��P�)H��85����0���^o4�ǀ� V��ܸOuK�h�P��N��Y�u��!K�%�ZI�=����x����R���{cu�2�� ȜWU�ǜ�b�c4�� _�U6	/�7F0i�����'֔�Y��H�g}&�4�iId�og�� eom��n���R�=�0̺9ڶ�Y�A�%b�.���4����M� ~K������廵T�P�Y��'1�N�O�ht���O��,�o�Ri��)�*l[2���b&π e�?��!�4\fĊTv{���<�2�+�R��X|xg.�չ��4�f�������u��p���B�&EgI���}��~���)9�p�����R�;_����	��? 3�.p�9\��@����l�2�'���
�����\�z\��ɉp�OoY��"d�h��I]�ޱUNy��DiC��8��Bu�>��e�mG��%�HK��É�L�Z�� N��y{�;�ET��%}p;ѻ0��Y��V�т;�����TB:|��k�>*�����.��h\���z�8&��sP�y@M���1�8�~��#�Ãi���{W�f�^�z��z���Yhe�=�ͬ���:7x��j`�A���v����	��L��Ȕ�<�(���%
hY��]���ڌa�Mel4O�qKe�g=pyF�Kf�M�����'7Ʉ���`=�E��� F�L��q��0=4.ǌ�Q��l�-9¸�~����jk�	%~���
�l�E���t��vDD�O����f�,�(w��^K����
4��Ρ��k-���>��J �]��Ic=����|�y�
�Ď�X&��9h�\�=�PԪmƯ���E��rKK�9�^N.�@��Q�2�2�"�J�r���ݳ����)�X4�;���=FVW&�X؟!�ಸ�g�[yt�O,�?y������l��2x�6�!d�� �rf��DV�
Rm����
 �@�-��Jezb88�I��$��K~bd*�����Ա�?iHsr&H>:�3�@1���ۑ��+�R��I �ۉ�VwbG}s/��,F�8��D��Gxfk&�vf'�!_��9?0L6(A��n����hþ��WRSy�B�%�v�ݺ�[�7�V8I ��a��Y���.�Qk\}#�wY��\4�2GWD�W���9-�p���E"1��ԓ������k�J��K
�8��FQ�/B���:�aH�PQfD�� t~n��)����R�+Q�d�{��5S�����2�(̕��"5�����ki�o�P���a��=���}n�e�V#���k�G�
��'�&��� I�×A���}'Q���?I��ܐgj�yC���jV����S�����4���Z�߈��r_�ߖg�=y4��N����A�|��{c��X�Nk�{�m)�}ot��@S�6+���J��\�{{k������C:��K��=��'X�{,GԀ*�&�Z�^���^��x��3�|� ����]ǁ?�j|�ΌC5`紟�l���'���-�f���'"Fr�ХJ��b�r?L�R��ܛl��?�x���n�T-5�|���h�JF2���`��:��B�}h�c��/*�]+dC6[E�A�?,�;�I��Xw�e!�꾣DeqY��K�Z}c3#�Ǵ;�k׽C�u�$��Ɍ50��C�����t��,����{�L�N��B��8�ޞ��7hg���a�>R=��i��pCWKzp&�|�$�̬�g'�w�\���H׼B| �xO7�Yy�*�����۹2��'��Z�է�9�q���k�!�6���~pHw|b!(�y�ի"�jǕ�1wc/rzTD�<Db��I˓�*�7�#��S�>������o��_OC
q�q���8�Of�⁬�(9dTd��=��������L�w	M��FN��Vhow��g�Wv>3jw���^�/��a:X�z�W�a+�2�]MYD��x�j�S�TT7T���x��(�&�u�B�A�������"��v���!�F˭�@��6/��t�bv�Ei�V)�(V�y����>YX0�b�y���t�i-S�A}Ʊ���Uj@���1?���_�d�YPU>��w�9v�����v�Əf��ߛ{�X
�ߥ�ִI�����mm���e�&�r��H�Gl�P�JUt���ʉq�ӄ3��K�j�Cj���0��{���-`c�TЦ��-��M_㱤&�O�g���!~��� �?�՗J���yl���;s@vN�<��*�Թ)	~��NU���c�����iB�N���R"�R'�'�_���}w�He���YLΪ�0on3�qM�}xQ��SϢ�@�dw�80�q��qR�hZ��Ź�֚з� Q̀�Ao���d(�i��Z���~奾_����?+�$�a�W���15K<��.h{���?^l&���c.}�[A%��y.o�ݫ�<�I�N��`���o]-�؃"���蔱�p�Ɛ�%����'P�Y�˂w6�k�ةs`rg�G����)]0�i�����J��.tR�b�Y�>�~͉���"'�J��-���b����4>�[�� �2����T�hi��B��W��[t!��N��X8)���h}U����nr*TT����xT�o������=����E�U���b�]�����jao���lq�
.�y��祺�͹(��E�0��Kq�n�jX���t-��E�"��w&�g�ye��R���`;b���*G�_���)�-��zKe?*�nࣂ��)t"~|�xfc۪��-�bI�F�de��a�J״y^���-���߉[yJ�tb��d��A��^�,����Eaе�[�((���Y�o�Ǖ����Ϳ��ԉSI�]H�>ޚe���p}�Z&n#�7����HA�R*$�N�b���"���2���FK��Ŗ��^�w!����Z:&�8?L5ޚ�i��#��} �d�����R�4�u��{�H9�D��KUJ8�{�]��m?\�-6Sjfh�v��R�=� Y�;���nL���-t�p�8Lww��wd�fb��3�r��^��3�H�O�����"�pMAIl�GS���\9*��q�ߣ<!�9jS��T��CF n�y=�L-��5+�	��l$�ޘ������N���b`tW�l��A`��ʯ�gG�ϯ��f������n��̹�aW���$�[��X;#4�V�!�5�E�b5��ЇB-���ab ���@z�>�'b�L&x��ǩ���~~��e�`*��3�cVa6���y�O�U?���I��������ޱ7��`���{"Sc�`�
����"ʛ��n��65�7����Q��m�$�ć���Ix9��K����#�?z���<�.������뛊')�!���Do��'bV۪��=o.�P���L�(B��Xb�]��P�K�Ȟ�E!OJ!@�:8X4K���
q{P�*>mp���/_�����'����NWz�v�R��/��"���+󿼟� ��4���.���to��d�Z��̖���ne,3��~�n~��7L�p�F��N��L���Y���|��ؑ�Z�ٙ����L�Jhg�Ú� "�B3���s8,�w�/�b�{T�uw�F��5O���-�O�o�JBp	M�P��$)�r����ƹ�]PhM]�W�q�"�ܟ�z�~�o��G+`�%12�A�U#�������%"޳3��C��ֹ�����W]����tC��	!9{�[��!:v���K,���|� ���6tP��A鰊!w��}]��дѸlzM�{�A)�e7�l��b�n��c�G�7��]�~��$��4����h��*fZ�7g��	��{�XTPc�P�cv
d�
�C,d]��7�BgN���;���@�u�x�'34FR�DN��(�>��G
�4<1�`�D�Kf������f��B�$G؟�>����k%q9]���������]8fj	�%:�@�	�%������~2�¥�R�o'� hg�_U6�۶hbvİG��le&8']�Pa?0G#t�d��<��@k��Y��0Y��W6�V�l�R��Vk�6]U�y�Ǔ�/7�m��?�~��wU�Ƿ���Y���تфxU�cg�f�sɧy�%Z�cɑ6���:RM��=�Zf���Ƚ���H �tjn�����Wػqϫo�6KP�:�5-Gh�9&��[�>#���IA�~�&�1˰%!K�P���L�9f��T[�,C+�V�T��~�YtHz(��~%^7��M.�4�2� ��n�����=*^RD�g2i;@G��Ũw��O��u=���MՎ���2�F�d|�"T�`ǳP6�������}i�r���ň֍<7�0H�7>�����&1��t�����n
����������ij�y�81~!ϼ�a�1���? ԃ�IG��g�����`�W���I������f)H;ɵ�}�:�w}e'/iV'n��F����+�ϓ�7LdٮC��ghJH��/S
��7�t�]���p�øᨶ�o�xO���-K��w�ev����@ JC��W�`�W�U'h���£�R�Y@!<)��y�]�-I��,��92O}x�<�4�<��"Zj��ݤ,kz�x���務�Y ��23�u�}���yGE��.r������Ԟi��|�c'��^�nB'Ҕa%�>7�V"=�'W��AL��0O�?@h���"4�F���flJ�7�D��7h7q�� &��jr.a<z�2�:4Q]�ϧ�C�:D�wX����smhL�Y�8�`ӫ�
(7��9���J�Z����v�sp�n��<ԕ����ɚ�������M�'�W�se�!�n�@�.0&�\h���35��������������]�E�) a���ڱ9�Ӯ��O�-�/���բv��쒲�~'�١�.���w��a���,���3�6,�����f�����/�T����2e��0�"�=w!�t=!�ґQbUڈ�
N�$9˒\��~>QQ�b6�$U����qUV�,p/�E��4B�Խ�ьVr��f����F��2�t	\�m� ʯcH�ɳ���9?;�]\�d苖��]T��$��Dn��{�!��L��R-Y�C
R�\����fP���#���!r}�}��V/�+H�x�&�.p���_7�� ?L���E7�Ņ�c�e�dw���� ����mݟ85�͠>�V��M�b�b�^�u_ȱ�J�W�r"���K����ȶHB�e���(���qzLb����m1�^"�����9����1ZWs�u���;7�i��i��P�!�wV�X)w�O/9r���+q(��!���peZ~�/֢��2��~K�q&���O�Y�!Q�L�\Ƀf��?��4K_�W}.T΋�W�)
xc.F⽬@d������jX:�K(�,�쎯D].�a)�@F�lLڜ�<OVLG��&+7��[��4�����N"��4�/T��y���g\���l������~��X��2BbG�DmC�q7�Ze �L���@�G��i����~�\�~Q��ni5zP��ռ$x����^�r�i�߅K�*��bM�6�=
�\�b5���N�1� ��z��!~n0q�����;�i�ym�Sא�Q%MH�}�o��1;.w� u�M`VS�	އ/($���)�n]"Ar؃]��[?�E�4��;��lڭL㸻v�l�h�x �F��'�˙Q���^��9���\�>'DlRo��r�th`��3��O{�1{ّ���	�^�FԳ�s�D�ⅇ���YEHJ%wOS�1v�"�JI^=�9[���w�0�_
&1���<�b���w���
���\F�n�q[;�c�܅1�y���?ƚ��$�ϙ��K����؇�JD�*݅=RN���A�J�e�.��y�1.��m�p�ꮆ��V�z6� 
�Tq�#�������ţ�Ry���t�*|XM�A9�}F����d^�/{/	��,�t�B��т���O�G�G�@$U �Q��� ��I�d�cy�	GHTt��sM�M�[�k��[n����+㳟��]y����`���<��}1��K�y��ͣ�#tȆ]�h��tTD��C�b���������_^��2�^���_���D�M���\�`Pc��$_�Ω��������[�?��������R�0�th� ����Fx�J1�f�V��>� �3�n�H�C� _�O'x抨��pbs�_V�?��R'J?rK6U=
;�%��S��y0M*��W�t��] ��Y%eu-���]�ӱ=�TB�YJ~��v%�-��<�N9�E�\�e��zGEI2h��Ym�ل�GW*�v��)��@�8m���i���d)0�~���V(�3������z��P��W6я�w��-Z�~ �GdR5M��іM���-zy7]��/�f.7���1U��wq#Lh����4<����xPX,uk7 ?Gk��R��!�c[�JP�]�L�3�H~!2��dY��l���%����(�Q����'O�IIl��Ɔ	���!_�.�Cb��d�\��Փ��h��X��-�Л>���=�m0]�vޓ2��	iN%���e�r�l���b�/�\�ZO�����D�r��PQ&�64t�8�����NE&�y>[�j���u�t��<Tk_n���|����U��԰�qJ�<I��I���X�	�� /��pl�t$A ٰ$P��G�qF�!q ��(W ��@$���YJ��K�d�]M<el�V"*P�qZv��Ư%ض}��n����o�Yzt&��7��5�X�X�.�c���ی������*��;�l�QN��ʮ`���E���:�%U�ɂ�:�Xin�u*D5��7��~<=�V��uًƻP���Ɯ=_F��R�t�t�+��(�<7&��~.�#�}|�� ���4kd�jo?(#̫��qd�YO-ҷ@��gc�mũ�jZ�p���y��H�9����mGX��+���^3cP�cd!��5 G2O�1m�ZF�:rX���+`�����J�z��$yvR����h�6kV4i���w���H>�9ȫ�g���r'=�c\jv�_����7����;��hS�/�_��S6o"���N;�<ʘ���a*g���Z΢��?H	h�j!^dN����%�e���PڸlcODR�@L旡���ǳ�ҩ�q�\��m/���p-HP/��o��:����j��m��C��rF���N3K�<\���lRar�jS�G����X>B��`��V}t��S�}�Nԭ����ңğ�*~�L��=C;�_���Զ��䖪B�h��D�6yԶP�`{�2C����~g7���}1º���q�(�n!u!]�v�_��p�!�A�����a����a/�%�O��2�c��lX�1R�/�)���S�}�_��h�H�%%�2�P����A�~����^|+;y���+d��]{����_6^8�/U]+���S�"�p��B�����3��y�8æ6�|5ǟ�k��n������8	����x?qtO�|�H7�
�_� ��`э�t��x�h���Ck� Þm�$�3�8n<���:�굡ғ�9?��C�LJ�>�������&�	��<D�R<���qD�@�Y/pN2|��I��̿K�I0�A,Ҋ�TN���;@�}_��W�tß\gM��9����ݤ�_7��C̚*�Ayf�w�n��?�h{�BRKhڂ@<�6bU����ǘ�|buM㵗\}U��T#�\�{��{Bf��@U�o�n����F_�=rq��O�U>DT�]��*��'/��Ef}4�-G��y��s-�%Nlu�S������]�T����l�q�/uj��L��հd�8��vfwc�v�֚/����v��Mi��y��2>����ѽ�s���~`�Θ^�
װ�H,�]�ZQM���y���y�d��h�I�	L�[ݾ0%a�?�F�)-!g��
`0 c����I����=��߫im�պ�;2}˷�>zc"ɚ���D g39���-"ư\�������C��e1����Z���k�i����"����X�'n��Qb�A�� 2��Di�7��j�FgA0L@��l̪�4����ɯ��$��-���.�v^zJZJ�I�AV` ��5�m�!��B��E�q�Jl�oȠ��2�&K��s�Ĕa����W��|�i�5�jO[�0(�p��[p�l!km#7-i�E��a~�K��A-�W�w�(�?`�!�/o	$H���Cྲ.���<*�L%xu���J��`ČJT������Qr�:Z
�;��n��o�|�\�Z�imE)���K}��H��0'����?I"�g�i�0E���[�-�q�6m�ou>�'-��I�Yo�#��v6t�r���d�8'��m��7�#��HK���iX�e���~ywg�aŌ�f�!�����Cc���� N�A�ح�[ ������W�Y�D|IսVO�˛w���lwHHq����$�\聤��*{dt'ju�HLr8���W�"$�2��`f5��Tʮ@�ċ4c�%	&M����3X�I�{X*i�M�{g�nʔ[7[̱��1đC�W8GUp�n�f�r�+F��!sg00j�4�@��T8�\�r��ƕ��$F�,\g��Q��=��BP�o�L�cJ��S�w ������f������iަ��N!$�=G�G
�UQI|������$F�D�	��h��:v�����x���- )d��F�[m(�zƨO�Xd4Es�U�HLWi^;�>~n!_zQl�Qī)���{��H��נ������0���
���<��<��_�Y�R |�YD�1�׾������k�\��T<h&DJ�����=p4REU}��C5%F��:ś݋�Z�E<��:�D��O��iP�U�U��P�=�}����;q��%7���-a+F���������3��=V_>l�։c���?�>���I\�n1��ʳY�����X��1�RC$
�ʛ���E�7,�a< ��UHd��qb�O��q���f�]YٍC�
j��Ĵ XW�-�_�C�ߠ˟�j��[�17����ү�F�h��_s����ǅ��I;tP�Rګ\�ݛV8�u��dn�Nq��I���6mt ��!V����!��n\i�]��Y�zh0i�nE�L��)�\c�:`�vCRXB�S��Q�Mb~ R`��?�p'M\e�ߒ&)�~T9�j�@`�X����:��eI7J�eSq��HV	oDh�Ϊ�k���9*�"L�3���nb��C�<��E>,f;��v ��~�ݻ�u�
_�aGe"�p�Ԛ�|�4��ߞc���+s,�,z��ہE�oο�1Ts�F���Ԓ�)�!��~6�]�Jx��>G�~�R0�qS�^-��sp�l(�GTRU�ﴪ+,e�c�A�Q4J�w�wx���T������&��i�jVr���9Oy��ē�z�F�nϬ7�.�{�G�"�F�j���	�`0�_ƖH�:j�J���a���1ĤBQ�����"U$��x��l^�\�Q��
+a�:K�{=���j�ÑP��{���>d�}ĵ��C��\5Y$M�c�0���a�����[��%A���{J,�D5���9�5r~V����l?�,�U{�Vf�nȘ]�_�G�_)�4��>{<�Ǜ��A-5�����i��w\�`�������J_b/����wU���c��̳H��4<Ƹ�C(7���^�������++�����j���Lj�d�}���}��kJ�XI�Y`�q���t�Enf1�Ak�ߜ�ה]U��	����x-$+��4������4����[�8�O��Lx�[CxZ\AZ����� H�.˟5l:,n�x#$h��'��t������9k�i�c�/���&;,�!�l�dά�?��`n"�V	��W�$�;IEk�o��)���\�h�|�D�`̳:����#�\�6�p��Nb6C8f�<�[�V��pa�t�lM��VI�Ĕ�z!Y��`�h�0�@+؞M�뎂��<|+>˦��L��DE�1��7��SO2۔�
Nf��O�ޞ�J٠���sp�&ꊘ���K�`"���l��v܊��0ib�06��=T��f�we�L�l���9V��ھ�>1�5���0w��'�ȫ���������F̢w)>�3(�޵�*�7w� Y���w}Yl�EE��.:������VI=7Z����Q��K��'t�e�C>x,\�E���F��Yf��i����wB�h֓��!Rt�1�*;��K�֐je�*���	1+�ĉ������z>AU�l.1����t����TOi1�h�ʪ�1��I7̋�B\'���6�G������ɔmЬZ��.�~�&ܢ���%�����3N(��~-1�n���D�q5/�f�̉��R9�kⵎ�0�������Whm��� ���}�5���|����Z�W���FU��dC��t:J�6$�t�\D*���\\��x\�<��I#"�DP����n<���'r���U���LuXkk���S	�e$��N:���7�<���3�3d��j��Ψ�1�M���L���T'��ݾ�#���NZ�]�Lrl����M����,�6����"�� �Ξ�wנd��|��Q���u�Qځjn�n�sLQ!�f+��=;��t��o��*��ϖ7[���9vQ�ג�]�t��{�F.��r(������,�ƳD������g�������H�s-VΟ!eWF-�k^��q��	a�YO��dp<���c�`�0��P
���I�z�L�*r?�9(K�9_�J�>�AH��B�����:h;<�y�/7h�-�C�����ާ�n��2��1�cw�n�Ă1�;�#��
Vi'q8�@�?~�C	���b9���P���<�Ƽ��Y}��@�X�Q �v��)3_[�y:�T���s��@2�BX�-r��H<1� e��&H�7�*@>#EBIZ��t%)�ĺ�#ǝ��	�tv�}�,��z'�V �6��$�ֲ�N�)�C�c N`��d��wWPC��.]���>�m;�rhZ"ώЬ�-`
�d����3�a���[:��6O���Y�7�B��|g~5����+G��ʼ}��^.��g��Ἷ��^�q|0IE���t���2�i�p��r�rb���m�l��o��}\�����#�v&	S�&�r�����t���ҡp\*Z)�b!��H�����Y,��W,b�*/p���Y\p��uZ��	N��pbL�`Qywn�A~��{�2�7��`<)AD�T�Ǩ��=�b���3�+Z�^���M���Jj�����?Yb'��>�U��m��F������=a�DEd���q#�t����(ɓ*q[B,��Ϗ���%ϓK��3@0Vjv�@1|:��o���"�Ⳡ�Ny�@qշ�5g�6���m�ܗS{�YJB�����]�w��I��?���',��F=�ǣ^���PL��G=�O	�v�ܫd��V2LUL�������5�s(Ժ^��t;9�T)C7:e�>�z� ��h�vt�Ke�8�i>������_(P&.7rw H�J&Ιh:fkz��Z`��͘��uv��g�x�MIm�����1�/��Rn��ؖ8��~��K>�^�#W��)�����ع��1L�>�v����\���f�r�G-7]�Ż���!���X|�֥�/�'�"��ZH	�S��o�P��[u����+8L*�Cf���}�뵓v�J֬-�ܿ�`n��^��ȹ���&�8��2���/������b}Qd�
�Px��;)��
*�������סL�2�`�\�]����N���x�F�pd��gZ�ya��\�9/��Bo�Ӿu[on܇}�^��x?�lF�~u6z�>u���:ڐ��MG��"��j�4ٍ��_�I���c�.�>��cq��3]N�.�!�o?��!-��fp�LÐ��@�1�)���t����%ɕ�b\�Ƀ<۱$���:�@; ;s��2T �&Rی�)��C雁�B]=�nu 8����Qf�1K ���%�K�^1Qc���z&����,�ֻ��	�Zcqp�01��aOG5�'�`�DV#�� 6��&�٠E?M0\���0�2��=F*	[���)����>-vX$�oj׎��� ���MW�dE����
�>?OY�����AεB%�t����0�i�n�*4&�]�(v�gFI��vI��G��x'��[p}��7�E�]��Mq'���?G�e�� k:���!�P��ʣ�� ���IC%8�oSd��\��C�͇N�]��g��F��8�n��'�����T�M����j$�r�֊P��ފTT_��1�2]�'��"���j�36X>�6c�# I��E��^>w�r���y���Q�| ���K���$�g�p�W�jd��8��\'5���~7���!u���K[4���Wg$5"�����2"��6���t�*2�������N#G#o��slYn�▉�7� k��Y)a�R�ϻ�_ۋ-R�0��K��ѐ����ɚ���$����D?����{��9�c����5�t�������C����g�_�
0���Rc �bn�m�72	�JI)C�j�©�>�;.�P���=S�f���3�=�D|���v���̈́u��>8��&nģ�`��{�ԉ����<��B�^1AR���k~�����=�?����]��īL:�u ��T� �駱)q$��im#����l��Xʉ,����bj�� a�8��(NH��IД���Y+�հ��_�[3tE��(gD΀1X5F�5�-Ҏk�ƮsK���Q�]@�� �:��:L�N tɴ�R�e"b�����|d>��LG�	�~�)`'�x�7����E2�����UaG�ߵJ�	�*���-�| �0+�$�N�����K"�7HN}N�^�L�������Eiqʢy���AK0�O�\8-:n�^�*�ӛ�w%�G抹ٰ r�؂Rr{z�!�=��z�����g�i�W@H���Φ���܏72��11�^$�΁?��QB٫��AB��J�h%W�3V��^B���Z��H5��k���m��fǦ.�,��ք�ܘƳ���b��-z��GR�H�D�oJ$ ��mG��tNtt#�
��I?*�{Ϸ�6�w#�m����l�ٚ&�G9̬�a-��U�H��Y[N��l(ݑ����4.�J��]�u]<M�\<kV�A��a�Bb2��Ӣ�yl�ĺ�K�1.�	��m�I����V��o���������K��	���u={�XNg�}yzgF�ՅWGGsp�^�2i>C�`&r$V�y̊��8�8E�vIf��i�6~AH�'O��0��^�\k��-�:d1�(�?������Yw�,HC%���?��gz�U��i�|�!�[�F�n�����Fy �@m�]J���8��V1����$vP<ٲ�3�&I�|�W;{U��}��?�Y�_?��^�Dw�R�O9��|^j�4;��4�rd��e��u*		\/�eZ��C���10'|�tS{f����ˏ�D�!���������D-rq��y1{I���vD���kĈD���:��؝C<u
+־3����ab4��D���v'��9�.>���N�ӕ@�Ֆ���$�iV\��2Kv�OԱx�^X{nL1�� ��J�hϯZ��ބcy�����-q�Y��$VF�$0)����(���<p�Vqo���T�JZsl���ɲ2�ۚqֳ4㸴���IS!qa��i�?�ϻ��ʯ���������,��~ؿ[�b����V��_�՚'cY�W=�$N��߷i5li�\�8��9`����tm����%{��$�Gv�U+��7P��eg���E�ի[�O �Ǜ�#I;锟\:8��.�86t^��ׇ6 <iS����?A���d�.Nk����
�#K�_z�˓�b�)a���*�T�ͦ� k/��%m]*�%��Oa��
�"S1�|���:.ثj�˙�qJ�����b�0��掔�n=W�^,������YI�k��O�=�af.'V�aL�j1a�}k(_l�{�����c�Ҭ��v!�Q_�7�b�w�/�Ө�i �D�J_7hY��E����(�`[���d{;�[���8��<v�I��kpQY�y:�O�su�3i�;�j�ʫé��#���*��Z�fka'R	��}~��7��K���y�W~�1,����w��}���0U�*Di!����7��������u.�x:���k`}��@���^u�  ��Gr�H�{n����6�Z�L"F ��9�� r{�M��1�F��p���Y� w�twl��s�V��/y��#�`m�EϠ��d�F�ެ�"�W4�,{+���]��S��u�0Po�UA�{���V-�q���̘��՗m6{�n��Is_(�`�DX
��ٹ��ė��<��rk)��c@� ����q�2�F�j��Y�ɜ�H�yf��c���	�������֪i9�VϽ��r����TK� L"5@������|ƭ�%�v�=�<�i���|*{io~��I�l�a�q�C���A�E� ��0��o����oL�+���3���`6�VF�(f��k��Uy�r�qͿy��P��nØ�Ev^��b�/�ĳ�?N�~��ĝ�5�'u���G�>[�U�4���� ��#jV��=
$�d`�L����'R�6��4m\�?��@����������X��O ����>�j?^A�����i	g5�wMQ��>'�E�F��^�2î l�-�	5"KYD��%��UN7(�(�j���4�L��e��kjÌo�9����#@�1\*�s�5ԥWч�RM����\�/��#���Ύ�'н�d��$�va�C�C��.*$�f��	��E@GCkک�ACOR�8r�B\���=����8�����/dL@j�ɦs��Sv����#Am��5 SPE��f�3�&_���#��$BoE_`�fG[���B�\��T���>���LM����)M����/و�"�(�ZTv�=�fr�n��QFv��}�e/�D�.�����I���G`0o�V2�0���!��� �G�|W�����i�ՙ=��O���&���w+wBE$�@nOC�<te��%�E�Ό�$�o����T'���!l�������/�͛+��A���ߍD�:m-:2T�����
���p_�-\hb��>J���m8�_xyɨ�N�ӴJ�M.�W�ַ�b����j}4��˅E�<��9�y�Q|3�`����˂k�\���>`H�2��Unrq:G�@η4V;g������3V#��V��?;�6�%��kB�ʢ5ԥ0�9�M�\<�)b2����7n�c�'f��w���$|C��M����GÒ;��@�����V��]��w�V!#�( �\F`� ���`	:�ߟ_�eu����N��	kl�?��z�<����Q��:x�r�e��e��������!M��KX%u}�'�>��o�S��4�j�
#����G�wi�jV	�0-*�J.�ޕ�5p\��?/���nz�p�*|x@G�U��L'�k��4O`��d{E%�Q���b'^�)�^1�Rg����^\�0�͍
4�g���ڼ�+m�6��3��Tg�ʩ��c���'s�Q�CUe�s����?4aX��Z��&R����	��0=�dL��{TXm���Y��:��h6Y�Z��o�˛�ө��_l��nS=#��Rk��P��N��O�k���c�nА��@�	�8C�{ZsxS3��r���}#�aP|61ީm��_5��G�%M��j�����r��-���O���N�x{L���ğXg%6�A��P�2b��������\��:ǘk
L�؅�`{9lA�,���ה�mm��)�=�,����'�x�M"��}=�i%ud��nMԬ���ޓ\��G��M�jf���(62	���|�d���K�%�(�����S� My��1x��,��9���TP���X�C��@p�����>���=+����rG�~]���j��VO�����5�I���Us��p
r�>|J�������vM��;�n���Q#�1X�%vm�(��|�}I� 8���@%P�8�>��*레���V!\�]��=n��Sn��w�����X�t���/3/��5ğ��5�Bلz�,�j���ppsr���B�q��o7��aE�xs��|��W���÷��J�:3���{�ΥB��j��]�~}�]���Hn�����<O����y�ɢ/h����!���P/���$�2f�gZ�������c�|�T/Iъ���;�uW*Z���?�WL[�H��%+(QZ[:v�*t�<�ؾ�?��G�To�si	'87�1�Puzq�>6�CQ,�!u ��C��o!�TUI����:ۑ�6T�XB{8�\���/2Eu��r=䙳�6��+�	*��k4�ً\cT��화��|��"ؑJ-\5��I�*�κ��T(�������MpU��k���>^�imO���(릾>t`&�|˝���\x���9��x7�K _��@�a�`�[n�m/��곥�U*6r�� ��qLջ˾� 䴽���^#�A���q0>w� �M�N��h�1?�",@X�0m��yM�����aw���i�(|d���k%��X�������z��C���\i�rڌ�p��*M�֜O%t?r�TGFMq�J��C�J7%�[A3���·s�:1M�*����g��վ����=�p���������G�^6��Nd3�(�~,�&l[I�N���������`�d��v��3�m�ʖF_&u&A.��Gݑ��D�11�C��-.B��64�$��
~����9l���ocᰞ\�ǟؘ�nam�8���F��3Q���@�̎Z��NM��M�=7aYU= �]"Һ�1��(�vGUT'M�s4�A>�,JyB�Wl.;�t%M�
�γ��|�9��S�@���7��������
��Gw��>��$g�S�m~Ì�?S�ܗr�� ��]7�1���Y��ԯw���b)@�3��C#��^ѓ�Oi�?�j���\��*�&��H���b6��g�~6��b+L+�?�� e�6�����%��Um�Ԝ-��^켏n5߿�_�@W5å�a�i��t�$��J�4�CćC$�-���R6�:�)\��&�Ƌ�� ��JO��/��l7�U@ 3Cj�Q�鸞:�"b�2��Sb��ꌀ�O�<V�B�S�?F3%�GU���y�!�W"���֘&X��4`m+��T[�p��D���Pϑ;a����=���E����*�"��bV&���$�tr����f��7��*q;��d"���A>�$�t�]V�p�gU����}P1ʳ���"�SULW��Ɖ}a���	8;���^`��̊�L �E�U AZ1��nES�`%�Z @���u�L���FV�-�in�m(Ӳ�~G��g7ZZ.���7��9;���DA��)D�q{��Bs9���?i$-/ǽ���nrν����N����gp�Ր��~LƔ���5������nw�U�`��i@��0����ט{���-;���*�sb��'������E<���4��H�ٿ�{+��5B|?/�dF���n�eEY��dzG���$;~|&_I�h���"�p�z�w}K)X~}Yd� ����F-�U�%����t��w����[���Ra[�*��b^�_��;u�%�es����r�yNd�W(�Og03n~��u4zd��F
����i���4���#[cF�3Ҩ���z���G���-�h2.>Њ�i (bb�	hF��i{�[�6r]"d��S���z��v��-яm�z�Ɛ�&��<��6t�A��)$��v&�'rw>o**8�PIs����P�@z4cR�՞Q���_x�r����J7��|G��K�HH�BP{j�dX!%�C�937��	v=|�J	�������/OKd�G���mi�|i���s��:�q���#�GV��ӹ;����:9�����$rT�t�}�(:��a2Eb���\�9�:;���|t�Vs��Zà�2_!���l"S���o�!Ș��M����cĶ~Z/f~�ˇ��5�D&�j��V{�š�c�$ߤb:���4({9�E7��C�za����\w"��#��4�� ��j��1���$c�hZ�]O}�eNZ���
���k3�ِWUw�*�bv��l&� f�3e��)S`����Y�$��/�E��u9����D-6/��������.�iTd;�$yCFE�a�Z���hW8��u;���*r����o5",D�P��9c�yT�(t@O��Zx��;}��� ���j���J��562�ʮ��Q��Z�q��Wwtc��ֹ�v"���]�o�`oiV]Z�C��։ݑϔ�Ru��K �fR<,/���Ҩ� ���[(���fa]�2*\�x��2!YgA;"@f�Q��`0Ҁ.2���������el����꓿���⣛T�U1F]�sFy�����a7Ѳ�䎅��Q�Pu2C�"��"��+�cd�d�I�Hwٞ��M�-ꋔ�������j��;�N���(x6[[�ڈ��M�79:gX�a��0��)�$ ���)�Եϧ�Q]��l.C`~����u�L��f��L��5�8�W��u�Ę	�- ������o���8Pfo1`JG�8�c7B����^L`!���tH%������B[_���m��^`e� 2&&�ݯ�J�����5�6l�ֽ�r"f�k��������{�+rWn/��s�b���c�s�:_x/k��j���U�=d�Y����42��g�\�	Y����c��v� D)�*���d��"Lw������
+�L��ӇY�q��>� ����g��%oK�f�ڶ[�΅��͹f�79�6����ۃ���+�5dr�ي�w��X3�b�,�+��/����� qX��ƅ�9Qu�b0Qy�%�'O̴��|��7�-K�Ej�\=��b98��-��?�?�)���6�ﲛ[�� �P@<�ҷmYXcF���ǝ@<���C�����
�`�"���q���f\0�D����*�)��uV���ْ%�W����`�ޙ����Hn9A��jN�A'�ڣ����--;$�Tf��k�E�G&�R�s�쨞O��7��7�c)@<p:���"��&��ɾ�H�����dj�&��;�.�ހ�gy��k�/���%�tfbWP�_o�%�]tI	z��[��膁]�=A`-nz f�Ovd�����ʦ� WLk�m�A�2�(��9����1������C���Y{��C���S�y��1;�w4���j�B��u�a�r��#��X@b1�?O�]c\){w�,`�Y\K��'eFZ�{#�	��|Z�
��0B`�pW@�[|�/h�7�ɑ_���}?U~������3�ƀ�H��v9�_9�!=4O%���ɪ +5���s"\S���7#B]��?�N�!>U�tX\�Z��%,�ؾ}bs�� J�s��A{�	"|���L�V�E
4��D��oY�NU�5]Y��?�q2V���UG��KmꟶH
�z�V�&m�����YZ�'���ܓ�$�J���*G荳����J��lv h��
��p��wX*}���(Ж�,e	0T�d�:�8 ���w�lh��舛���G�Oψ2^�|��T�Iz�IlԵ�ɥ��e_�c!��5빫Y��uw���"w�^-+$�5[Y�5�"�Z��iS��w�YV��(c�$��]��v)��XC�%84�?ʎ�BO����^/=�|`Ǫ�a�3��"ZP!l��e���6�׎�n ъsG�)����#oTBu8Y}W���!�2���D�ޛ�Ժo�5�o�:o���:�j�GUZ�T�{ �������#'��B�B�$�~��,W�
L��zy�	{/���8_�]���'�Y��;�A�Ks�B>�t�#���$��,Q>�21ǽ����5��O[&ԁC۟��W��	�hr)9I���˸�2���|YDV��͢�CE��X&�����dP�]��c\��'�Y�v�灲���|�ei��m<: oC�rQ�L��)�����:D�b7��<-�-�����ц�"�UJʫWy�z��^��M# ���6�e�;� �>ЫM�e���}���R����S#�,�l �� �9��Yb�[�ș�vԟ]*3���&QN�����t�?$�Ɇ2�G�U�݋*��0�A�+��*K|��@"�E�ފjMU(�b�3��{���{���_D��_y7
��@_��<�V�W����=L��wN��z"H��\��x%�?у(��T��|���s����U�qE6�>���sM�k��G�� �c��Z�l"��!.;|��R[�eB�Sd����[0��t"�P;`Te�ld~�B!���
1�٫�Ӟ�D��H\-Y(閒�*�	�����1����o/el�r��j����]w�
R�P*_R��KzW"B�X�6�5-��Ϸ����z2��-2<j�P������jS��a���v�AN��̽5O�:ѽ����
�7�?fA������2SU,Q��<�ڈ��8�U��>��R��w����S�é�4[�q�n�R��\��N����� F�P?�������k��eb�7�����}�9X�!BM7�-��l[�Ю�4(a�{QUXh�#ťEV|&$�^y��Y6^���P�X#L~7�8p���?�j\�9��i�H�(�����"�yf�!�Y������-��<����:��L�Cq.#����?\�&�ym}���*0m�V�#��y×�W6Q�W��l����s3�ʎ�h�X�@����K��h^�¢b5;��,m�i���#�	�tl����eVQ��t@�rkbD&d���wX04�`�����y_ִEw@�USv����o%�q����r��t��4`GT���t�ߓxry'X�zX����X�oc,��[�����������H�!/�0̖JT� {��.鏥��k�z�4���Q��HA�m;;�L��������5n4�8���.�)o��� ���85Q�9gh&gal�??����]������ �����VLQE%�X���bH��;,��b�~�q�Ƚ(Y�ܒ<#�֨t��8�Q�a��d��Y��ϡnzI��|tN.V���o/�G�3�w&�8��+�\���%8S��_�mX%-�ڒ�c�Co����0��
�<���:]��H�63�����I��p���Es����>Wr ��x<�{.Q�T�(��z���s�?��.�%����f!���8v^���k[*��;]w���i;b���,������\��'�W� k�H<�q[� ��Ɇ� ��3�rqv2�eڗ~�m4ۨe�9{��^����p�	'4�X�<�Ц<t�sx�.���x���-�E��ZR�ҧUvQ�t�ݴH)��Eb�b�HR�F���u�_vBee���f`���`������[�֢���x�:�C0qvu���~��)b/����=�a5��d�?�s��o1ߺ���Ј�Y��8���QS���L��j��gw�pO0T:a�=�F�FYhd�ۚ=̈]��7����(yu��w0Z�]cK\�Y$3{��螫��ftJ���燯9��ǏZyRW�����׀�HZ�k�A�3��!P����������.�u���\!�ڤH�����i��Vk����t������J�ŗ��)V��mﴻ�	�_/���aI���y��Ui6cj +)�E#�!����튞�-��|�z��N�Z/�����~��&ef%��^S7�ndŎ��-�\=c>���H��'iya찖>h�����Щ�;y��4����ZĿP���N:ݥ��Jl2������W��{#��%S�E_n�Ba�-h��E�����@���M� ��d>��23�Q?M�#��J�3�Ǿ8��h�_;�6�:*��b�Ъ�n�y�-p:��o]1�,-��5��ۊ����X܋Z�<A��Mcp��y�WwOy��{8S��=���a�G3������7]zeP��!�5�A8�^��%2D����P�>[���������8�M+D��˒�}n@�
:��^�X�_���T(�vB#�I�[|Y
����+�~v��T�
��M���lɖP���v���x���
����,jq����0��3�"�l>'Wʡ$¬�Ѥ9���;�ꦛQ���������������K��6�����c� �N�
t��I6 #�/BIAb��"sr�U�n[��Ke����bW`|�Z�9���8�a�L��\7F�f�ӳ]�C+�&�ΖPk| �9�P?�7Ȁl�>k�Zb��y8�=ኧ�����T��F/�x�
�j���ם%M�J�\��$�닮g)P��De� �u��������i�k^��Pe�U}D���R�ػ"��	�d�C �W-�*<4�Q���	T�,ށ���:����S:Y�RУ���$-��*Zo.2�#�Ιq֪�s�)�v�<�UMyn��xŐ�	y�¶e���N]�A��!�mP`'�'t�a����X�=��]U�;@R���'�����"�6.����Vӆ0�r"��]��S.S\�q�I�~��ܴͽ��ެp�xBڕ��|~��T �/R��}�pG.f���/:��ӟ�7��	�o/��������)��fY�.Kai=���{����h��.0�y���@w[�E(Cƴr���W!C�x�i��1D���RrSx�s�fYCO��Ahc��g�&�;�c5���MI�+�v~�� ���Ӣ�[��c�F���:��onHw�+�QFJ@�{���0$K��'Ņ����,�ܗm�e8b�����0}Z���v_�g|]�ò�8G'��m�NJ�����t�^p-��2���J����i����}7�Rk�j�z���&�}�(2pQsf����)R^���Z�(��L�pM��[��YǑ�yqDkf��l�Rǌ��!����	7��(���خ��j鹎�A9��Ò7ύ9��S�&��F�ճ�b��$�-U�ȫr��K��&�F�U/�4�sX"C+�A6,Gg�8j���!����#B��с�ә3)�i
J��	h����3Ԝ��q�#���/�O�\�.�o�J�Mź1�xZ+0�ԧ�ؚ����F?��1j�Q�\;xpn�;�b�����(8����#r�8ݤ{W3=E�ip:	��7h%r�Sp����av��ߺ.�?_�0 �_�z�)��}�M����L�0�޶�(p��)�i+�k���Aj9���wW���3VÊ杍́l6����n�W�+�'S���T�9���]!���Jz|���q�ѴB,�WB�o
�l1d�v:�!+���,���*r��p�����V|�fUk+����J� �-���sw��۔��w ���*�b�Yg"!�|�}
�G?o�҈u�
��y��G�94��0�Yf~���9��g��[�^?����΍%���3������~�f��ETv�R��a�vϾ	ү�✸����ͨ�)�t�<+��c�����g���n����*"8k_{>-$�d�{31���@1�ұ)k�6Z4O�3��qvT��P0N�C�c<�u�Sd��]%���^��r%]%�fb3�hd���m�1�IX�}���!n%g3�#��JD�}�ޒ�X�e�q��A��4���>�QAL��ۍ��ZՊc��'K� ������m�������;?�,S��e��J�Р>��g�#�q�\�)�,P���C�>ipQ�|��2�y@#�o��sB�U�#W���cuUۅ��}�q���4�x��
��dw+o�M���@��5yZϷ�S���l����XSk�cҗ��
���S������e)��Ѡ| ���ԓQ0Te� G�N#�VU�p��1��Zy���v!��������p�c_��.����4%Vc��!�p)ˑp?���C{1��@�[�����!�Q����Ϩi��\wM(��3�nZ���6BU˶,���4�����E�{�*]��r
3s;�4p�:��Qpm0�Ɇ����I�vz4{��%ZZ��� ���7Q.0]��&!��=k/�!k��}��jOK~�
7Hᇄ!�"������:j"��-��7�P�"T��Cq���Z����׆ ��r�2������`o����24si�1օV��n�q��{���{ӿ����b=V&eVTq䥩L�1�_<ʴq�؆�?g��I-6�!������U8K�$���=`L�J!�k��ѵT!_�֧w�:)B�Ѫ������<��r~�\ �<#���Ɋ�_ZY�Rpii�[z���1�Z�x�^�Z�x�V�Y�'+M��,�R�E0`L�N(��+�/�o.�i1�Џ��������Q�x�0|������~����޹�! 
�O6el�hgP_3QZ#��8s �Y��R��\*r����pź\�mH7[��`v���a�O�w�c��� �%O�T ���A��z��9�^�4!'�7����lFB"�5v
I��.��"C��8�ք��߫�(i�1���c�C�݂i�璗�`Y7m�=U��86�>�6��;��P"�����Pz����Y���ɹK'E�����om�?h6��N�o#>����6cq�<�yG8A����v�ν��$:���D����hE�'V�?���8Xs�%�±ڧ������4 uũ'b�z�_�,vĕ���M#E����Vf�p��/��dd>2�ķU(���9u�H�����k���x?Q}B���]���8 �(�Leq���8!E��Y���X��ίu���%�����)���x�rC���[�,w:�@z଒Q��)����0��j% 
1�	A-7�?R�����@�
��as�1�q*W��[;i���ѹ�d��v)���Z�|T���,������-�Vp�UD|�(R0��n��k�[�M5d�9���� ���8��l���9!��`����K�ԍ�,�P5'����X	Rwx'���V	wi�59<2�bW��6Z�[����>B()�N�H�0�S�:�A�S�1�%��^��͊����V�U�+d���C������A~d����NAR3�I�@�Y��3q��f���g]#}>|����'m,�4���X}LY.,h�_�M��<��m�s���
%�"���?)�s�\�O[@���bߏɛBR;��>g��9�~���!���C��C��4�)���l�Ϸ/��#؝��7	锓ej�n���u0�>�M2��aj���r������nO�¨XN�y�?�bMuJ���S.�b��X�Zӂ��L����[<��&�/p�=�=n����z�R�<��`J�.P�V�#>�m����=F��*��*J���F!#���V]��J6�E�����;E��� 4`�{Y��� 3Ƭ2J�@��ෞx�#������V�A��|O3��<���� ^>�ʢ�,ʹ{�IT�Q�ɗ��z�oIf�� �ٝh��|�W!Y��5h�Ӎ���~��a�����"b/���W��8�9D��Z�Ȍ����e�����x�Ȣ��KkA�m�,��<%6��U�mk�5~���\��`C͚ƪ��_�B�m�c݈�KX��G'W"I�@��l�xQ$��ԍ���1	�H
MC9�yrb��V8"�BaK�c��톢����R�R�28Y5����oߏ�l�RV5~�&"g>q�<�t�w�7�[�^;��_4R�z�z�Lq��MG�#����̬��y_��!(keɠ����)�(��N�����6�)8u�	�
	�DB�\t��D��I�.]���s�
C��~b�:_�i{.[dVU�jVLb��qI�����G�*����Y�m���D��>�K�;�TӦ��OT�+`�|�s�h��uVd�vH��lƫ���#[�[�wa=6˯)�uT4td�Jnm��v7 �W_ʺ���{�}��<ѩk��z!��<��L��^�M�i3k^J�#��&����;c��V\�O�{�2��� !�����Q���K�+�.�v������J�A7Wu{�Iw�o��_���s/��̮�bN;���?������Ni哑�G�]�N{t!��^ۯ���A��#��a�� a�S
��ȬR��u�-:YQ��a�0�愴J�������i�^����n�������T|�K��dQ�zV|��Y��~m}l>���\��j
RX,��0�*�EzA֣�c�`������)̺w*SA����� �hKK��b����݁���U0#��"R�QJ'���UV���?ɠG��q�I��D�������\��C ,Z�Ms�Z��E�q�2|���(e���܊��@��H~�K6hV-̣xG���{�#��y�4 Q�[�+�x��<��8c�-�(|����OA��|���w�')��	]R���?�۾~_A�!��rҹ��ls);?�QO�1�vӶG��
�ߎ�eW�#��x�d�e�h4�1�i�m֧��8_���=5/k��[+��'�.H���nh �5��\���O�}�R���Tz��G�]�d^���P�2�c>;ٿ���ڞ�b!gA1q}�3��A�A$��A���
P<�ò�i��d)��wBs����%��.�	����4GʝM�8� �%�cc��,KP�3�=Ich f]T;���B݈���+{U{PZ1h���gϤ"���O6.=TM��0�멈���E^ ����8^��a��s�Zv���ZS�gƦ�U����V�XH�!2_'`2R	���iS���R2P;_T����>v�)�n<u"�U>�ô����4��/Igf<1=dY��)$}�z�۾�K�����B�2<�oܜP!��,ȄE���B,�Q̛<�]Qq�V�^�F��/��7�fپ Ѳ�M/��;�}����C�u	e��ީ����}!J�D�
h-�ڣ8cB����R�j륦�|�1WJ ���3�%H�Ļ��X��b�%�� �Z\>I6��T`嚍����ķ��l[de0΢�^n|����Q\o�d6<}oN���z2ݏ��Q�1��ԣ���Ne�\���Z
>�aQ�B�B?%z�=SG��:J�W_��7eK,@g�����~o���"���4�Ig���\�w�}�J��e�PԸ*�R|�;O($R[���Ef�NH7х�y�7�a.�+��g�Ll4���5�1����+/���?$�"�1/QW���r
7�/�1�|{=��A�mR�N#l���]F<��)Ǫ��(|�j"��T�l�c�K�o�2��(/'E���4?�K�A���Ƨ���s���A�p!�QAB_u*���vK=N�4�Z�����d=��1�+r�0o�y'��KB�N;����9�7?��]��t>�8�}E�t���֌�6�5����Ǖ-Z�hW���:�쉊�+2)r3��0��ˌ�YL�X⊓Ǒ8�\۽�_o�8	|��qr7�j�Ϧ-�JD�&�ѐT'd���l�D�J~�w܇ 6�&�e�3����K4ѷ�����s����;7(�3��\�m����v�G�[]�\v�A�y� ���+o4�M�ϑ7cf	@�f"�?b�i�h��nh�W���y�8R�ʯ"�Ğ�g%�J�� �N⠖M�9I�����L�	���%`xӠ�b�P�E�,��M ��2�L�J�rCtW>jA�H��F�X����1�6�*A���Ц�Kh���0����K!��-��V:n��
�\T�����w�ɘ�G�����vo'���G����i�G��"�׷�)�ë�f8e��B��Ԑ����:z��g��6�R;�ZK�M��UuE:XFpY��3�<t�2�tpɧ�EZ�q=��>����P�z]:Zu�l�����	ŕ����/�2�eŧf��ӛ6 ư�,�L�w~�& �����W��D�j��4KŬ'^����@f���z��v���o�5-�/�=����[������83��(�݄�q�� �%�>�y/�r���G���c���bZSd����­������e)$�Y,��z�a��x�Ųѷ�����]�����޳��I�^Č4��Իv�5in�@Xa#"/K6hA�q�PU4�3V��g��ݵ�斵�ۡd;�v���.$���0ut�����[eD��n�r"@鸞��b&�?�U9
�%����A���&����}_�z bZ\����/�,)YQ��&D�i�FK��!����,N���}�e�c,F�e1q�4u~�/\���?o*�أ�(�2��dӄ!�F��
�xJ`��=�y�W�G�x|������Us�bB[�_`	`��;k��0�{_�F�r6�hS1��A�2�����T�U��a�!���h.wΖF@���=)#_N�3+?��a��u��q�����"Sj�������ݟU��#�j��#�5a����à3����F��W�Bc$Dvt�M��J�*�|I���-���V\���D,A�C�"��#��-n �l�Z
e���A �8�� �t=\��9��V�]�0,UU������ �9�u㭔�*����s�<8`�����1��N��i>�)O(��X������O�϶�����󍲝d�B����3�dB}�v�Rl���Sv@�0f��GiX
S<y}ŭݙx��o�+v�;QV��ʙ����	�˫Xޕ��
�Hm��4?�#��y�QG'�#�v���5p��H����U���/�I�@��B��YU��W`�0�t(��ͤ69Ł~��rpk�ǜ���"~�<�G_(#MM!�(���_'D�$
�H)+lz�7���'��
=���1��-�Bi�0�c=���InF��`/߱�t����r��~.��n���~�FZ}�=��~u +A�^$x���F��R�8-^3�~��`��&%��@K�Y�!�,�6ϻ���g=��['� �7/�s�9U�Q�6p�mI�+��G���̊�CJa*�A.�{z���$\�d��q��/c�i*I�_Qi{���$47ί���Q�MA����8�E �Y����{!��1p.�Ѧ��6ސ���H��.j���Z�e���?��xe�x;?��&�h�d2�h� � /��Q	9�Ϧ�r�(I{�IF\�[5eu�j����q;%"���0�!����]^�4d�
[љy�'�x�Uh�=�(M�{(멡�J�'�`�2у��Hc��GŰ�Y�d�����_w�)_�K���5H�cpx�u� ��Ά^�	
��h��:��P�=�Q�$�r򰤻UkЦ9U��I��CZ48n��z;��E��˒�Z��|M8��ZsAi�~�bO\�{��u��rB�r��3�'��G�,)fje��n8�l�jY�+�x�R0�u��#�9f'4#_�S4魥��S2�PyX���Un�Φ�
�t2:r�$.7]JVVSt#+�ȖD:��b��*V�S�������\�GH{]�,�1W�r:D|	�}���,����� ��#�c�h�d�Kx�V ~�v�5�Rz.]���U��*�o=�����5ZVrr���$0M��k�&@v�.��4�ȩJc:��P����@�k؁{#y�<���}����*�͸أv�4�	��FhL���30A�o>�W���:�9N�i���Z� �:��+��]2j��RH5��/z�����r�_�%P�ġ�0��~���o�ڭRρL+�t������J�����h�Qے���	��=#��ϲ�'Ǐc�V49u� ��Z�	!!��������n�����l�ŵ�������m�'�҅*���6D��&W��Un�pO�7)������<����FZm�4��GF�u����3v�r�JQ��N��^�� uKzR!G����vǋ����
W��e���-�#�7Ԯ�)�M@�P�߬5��( wͼe�����l���<t��Z�N�9���i<	>u�)o�p�c���@u�T�0%����D/ͺ�=Q\�1)l��,��zóԻh�<Q~���!����YQ�F䨏#M�lwM�@�S:m�q�M�Ķ�7��`1q!S��Уj���2����y� �qg���isW]}ߋ�6��7��7����m��#��O���+��J����
�	���H>��#%��k��)}��C7;��p=ц@���H��T�Hr��De��n/�p�,��Q�$���#���YgB��"�En�%}�H�%���쥫��T'�/��'��,(R��e�]�����`(EK�W@�4
uV����S��û."]���HȢh��K�Rn�ngF����7?�Ć
{s�Z�ݲSV|���}�t�qf���J�Y2�
�t���f��w�ev�˻�詟�m����6"�0�O����z�t�S��7M�5�.���RK����dY��L�$@bq8% \^�^{�E�g1��&�g^�Ĺ^��� f����?o��t���ҷ3{HU\���`�y����+~���� ��Z>���V��g�obh����lq�Io[r9�N!��T�%��[k������yp3�P�@�n����l5���q����KQ	�*�4��Y՝X+�F����W�K�{Ѳ�)����!�g��C6�P �ͣ�8L�����z[����������}W���T-�=Ҿ����D\�38c����9Zp����
{P�Q l]<�K{el��ᡮ�G�"�7�;��H5�$��*h"L�G�Ri�����<��T��:�&T�)Ȭz��,����!�ri":ť��G��z�$.9�53[�)�OF�����ݕ1y"3�F��b�~����3'$��\ �礙�g�,�s���+�t������z��<�WTM������E����B�=P�d�� cD7`(S~NC���Q���8�Yh��˝�������5c�¤��ɝl��a�/�}�P* ��ht�iK�v|�'�w��;���gJT-f�M���_��&��DbDC�������pq�F���cAy�0Ei3_�G͓x�*߿[k�4�p?q��苒�P喖���8��m7b��~^�!j��?�-`��2��ֿF�1��/��	V3�S����>*����^�-?���e���{Y	��sN|�'�sp������)^�o��̦a��Q�m�[����>W=��[�(�P���jH&,S�!7�Wqd���p��y#&�x/����qu���3"�T{,�
��9҆�$�����PPN(�le�Ul��v�W��)�]�-�����>��K�xo6~����W��.��W[ɢѱ���;[�75�t5��&{E�
���gI�i�03���:r:\vm��IzHk~e�G�I@��~�/,���㡊��X�p�:�BJyj�w�\5Ͽ<,�ې�˄~��a!���r�&����lX����a%����/?��l��]'�yY!�9 �[>E����G��q���|���*;Z4�
	��?!��;$��e�JVi�Y���0iP�E�?�YPe��,�l^��3�q��烁G�w����b#�Ϥ�W��v�����ӎ秬(�m�)��"����Z����ڨ��g��T{/�ݕ�P���8M˿��/G�9�h� �D��_�.�8BF6rz��D J�V�: Á�R����	G=�}��
��L�&�Hd�����?|�"q	ި����ew(������2&z�a�3ځ0@��F�[��.n�
!ۣZZ������"���cyr#�X�&^�����Z��q���4��y�x�2dIB�ݫX�#��~N����Lk��cT=���h3���"����Q���rH��`���5K��+(�I^d7��ƣ9楴wE�]eL7LE��]��MZ<ce�o��>����F�4VC3GTՓ�x�b
��uVZҸ�i�Z �k;����-�l� ~��+�梼�����9B�:p���LO�ɑ�~~W�_�EH��~���dM�W6r�[޳�P>=Ot�B�g���h����,���n|v�asMaA�Fh���(n��N9ඡ��e�U���dj����[�*��I�$C�! �m쭻��f}��,zS�H���[doD��j,5�N6��2���F!���s�G���e¬FPWҔ�T8�Iz �z��pV�3r]�u{����_�Eu�� q��������`�d5������leC�:��4J!˛��qq7�H�وyZv�p�~8���;ً!��Ra�x:=\}�t��d1(W��B~q������q��A�§���8]��#�HU����\�/m�o�*�?�$'���x]��@�u��'�=6�}M�|f�l�.<���k �vڐ�W������5zU�p �#S�^���1c
��e��,nR%�c8Α�Q�f�W�Y�⛑�)y��l�W�
���/:MF��N�c��Qf�Fsl�0cai����������lg�1��Cդם�JVz�7�!/��gG��a؃�r0)]�=�ʛSJ�r�%ϐ��yv3�U%W���m*��1��h>��wS��=�����[��������Ca�%�QW�Q�1�����F����S���py��\�T��AG��G�,Ԟ��ފ�wW[#��L�ZI۱̹U����1����n̲�P<�M���I$iᯥ�Shխ�tnz�(#O�$�z�:!a�8��J��Ӎ�8������$��g����h�I��jvm�x�J�<ː���9���r�)������|,��vZ��v80�~c�78�j�0�g��/d��_z2�I�%�ח���5���g�J����I� q�m�����v�9fU˱ )�9#�+J��v 1��G��g���@O/���ϸ�7�4f m�%gJ�,"�Fua��|TafL �\(���D$OH��sԶ����灊[y�U�{�{8ʳ��k�Њ�*��Ob�j�~��D��'G�>���s��^�>F`3kŬ�����}�_�t6�و�����a������o��h�&�Ae8��+�sa�p���B9������1����M���wO�B�;���C/�Ñ8�n�dJ�VK���U2_�6�&D$Ú�d��b�x5d��Ιw���/�`5X/p��J�&� ��gDcC��J��<��̗���<I�8R��6�3�ڊ���Ӳ�%���v��F���VrQw�����1%p���|�3�޳��h�|vӉ�~��G��j��(�y�$��~�5�X^ag�u@�U�=��*��<@1�}Yqh��=3K�ָ���}�E;�*�t��s��d����W��N��$�K�=�����X��2�Z��b�n�
�E��P�4�Q���9�˔:']�n���yW+�J~�I���2u������x���mZ�G���`�i�(�3Kj�GO"����`~0+��@N
m���4H�6�� �̓�b���?����n�m	A�M�_��Cɺ�8�ޙ����~�����K@N|�Y7_��%ie[m�$�6�q;	04����<�'��肎nG�o�$g �3�#�B<���F��xV?�������hXOB.|�S¯?����H��iK~\��eۨkf��2|�$��T���W�L5O�wE=eW�T����5U�U	�V�aI+�O�Qi15������E>���`�x+�qHaJ���OH�2౥	>Vz_���k�X��^	�昱!ڦ@�-_�(|��)������h�4tB1?���[��[��[B���q���z�8h�p=e���A�=���^��)f�����>|��F����f���ʃ0��ιV��~��#�:��M�G�vYX�2��(��W��[V��L�o d���K��QS±'��ڜ�VԎ	"X��^6��gY��SϢ>�n%\���RI�itAw���� ��H�3t5��1𹯆�w�%1lg�I=
;.�m�z��<8"�B�$Ok�ǳj	���?,��I�V�S ,�%�f�Qe.q%�Ě sz!HQ2ïj��ɦY�Ӹ˲�s�C �^���FJ��po���A	4�$]��G\��8B�Iя���qp]у\P�?��g���I�XaA��A����~�"�_�J���RR|����?���<�Y�ْF��fCX��-x�z����l_�
����̒m?�^���*�(���&�"E��r*�c���{�dB�;YS�2��=���H�
���I�M�E~�i$��֑=R��u���3�G=��R	Ǘ�%$W���'/���"1�*/Xz��%?77��C��,^�0Ň�Q�5�G.�?�\���8��&`�B���S�U��c�޻�lpDÅ˪�<_�͐�i-��B���r3�6�g9vA�C�Q'� �#"n�rR}���Ԍ�.Z����j+�n��oC���Uߞ�I��p�]�J�x���q�i�*�՟��
���TBT��d0�H�4(�:ǋV�l�����'���`��5�g�G��B�j9L;�{I6�9� �hx�N�ꁞ���(��h��KVM������P|sx�G���{�^'ь��!S�ͦ�;A/L%'`u����.�Qޮ�M��l0�O�8��JTR�y����#� !��q�]�� �g�ԏ�����O�E����cE�F�Xlv�kk��a*'Y��0K��0�n,��Z��l'B�n;��vz��W��HH�HП�T�s��ĝ�+��i��swb�S/v:����>�l[��
���n<���L�?�֧��T�I�t�����P�O.��az<��BB>�.pˈ\����[���0��Ǌ�
s�.�2a>^c���Q) $��K�m���w��#��J��/�ɧ{�>��̒`|m��ӎ���66�4]�����D�KQ�S�=�g�oX�9���$U�p�r��kA@����5z�N��ʄ��pjX�'�F���}j����$�U'���-�?�%
��BH���$8d����YX�ϛ�	��#�׋,�4�16��E�o��yR���Ҿel�)X�r���/(	�Q���uiNX��W������[@ax�Zr�V? �d���1[��c�&�2�0 ��YA.a������bϜ9���A$�몮�.��O�� ޮs�곑�a%͞>[���[C8�8C7�i������@1t���)� 'F�Ȅ��������i@~�,M�폙�����`[�+�U#w�p[H,���<yd����sw ���>@c) ��7c�I�\�K�𴌢����MHJ���v"lM��0~T��2��.` ��{F���SL�<X�NW��/+����Ԑ��bL�|:Y>T��'�����[��H��u˧l�t@ �J�s4�Q]��π�a"㩽cM}�.3@��6Q�С�5$�lAM��V��y>��sD���df�m��ۯd�l�B�#PQS�'�O�'����x�´��1�a2�f#��)/;H�1��H���5�a�Od��Qd��h��b�����N�5U�(��:(+��Z"�[�.m�jj/(���F�ɤ�$_��bb�#/}�2~��x�K'�4�8�?s�ܓ|ݵے��߳R�(g�k%Ir��ŀ��t?A!r
�������U-�'=�8��|���G0�ad��=�ҙ�=���	r�����K�Y�8��S�W�DR+�]P���'Й}�S�>�W��+��v���O��/v�̀	�T9���h3�3�O�H��#��
�טdGkV�ӵ�F��o�ɹ�M[���Z��U�!w�찜b�;�U�)2�(�&��R�B�9V@��l1���	El�Z���ׄ�^�" �L����e�h��׭�IN_����c���'�R�ǽ����#2��ȷ=^��
W����k5����@���;��������FU'��6v���I^����h+:��B�q�Ǩ��"�M���&��yԃ!�!	s�.�s����u��=)��y�t����yI����x�$�ߔ��w����-�y$�q�W�S�(
�h���K�j㴩��n�i�����^H��ȶf8�9�5@h>%r,�
p��q	�Gm���,� e<�!��ܳ��Yq�ZymWd��@`X��Y؛$A��&��n�׾jj�=���X�38e��M�rYLF�Yf���0m ��8�5�G��Ro��GY��L~t>�W�Q����	 \݅��3��b�`�g����-����ck�Bg��G� %�d]�.�0�L~o�&���uazdP9�z	OmZ�xI6�1D�S6M�>�R9�Eޟ�����-�4��!�W~���>篯sl��~�=Z���ҲcD'�ą�̥��w +���on���gQ_��訰ZLg,���T;��x�pڊW���}�$D�e��uؖ���4�.6����35!d:w�m�%���@Ⱦ��ջ����=(�p��o�ѧ��!U,�L���8{������\��ʽ����utvF��Yt^��0%(��;�����WG ���MuM��;�(�BY�[�8�~4s1n���}�H����l#�(�],V�V�:֟����藹Hi�Ѹ/��;_�*Or���Ipt�	ç�9(��\w��E:�]���d`g��(|yVڦ���d����t����/y��c�!Z4a�_����LX��R=`v��ѣ%��p�3�;@ngݭ�������0
ϒ�m%lC1�a
$���$��ׅ��[ʝztթ�.i��������b����Ά��"Y���&aDD��g�t���f�+�T1�^Hc�P�n���_ڜ���z�Z�G�r{w�r/Ӻ�qGv�C촆f2�S6�Ա�v�c%���Mv�G�*���$]��sY����n(�-�F�/۔IkQbV�u��=���o+�5^���[�������Uvf'�cu��\�',~l9�y۝����ƁH�jjԡ~>��w?Z�q��YIT+�8�)��)��F�~#�q9h]S�A��+&� �.GV�x����Uf�V ��ʦo8��UCP	4�����~P��S �PL���*y�����L��������K1jnݗa��R�ա��Y�Tc�<�4П���1��_��^y�\�rdC�C���Q&՟y���\,�=kۖM>Y9ޣl ���r��1�����ҽ�"S�>Dsx��?l;�7B�������R�59�� ���1\�1�َ�������49U��d���|�wt�E�p�[<+��)�$�o����>��ȸ�r�t� �
	B�3pUw�)%4�¯���2=�D�Tr'�s�S�䳞]��(�v640z�����m����6���%��3��//�3�N=�p)!�B/��Op���rab�7����t~��,"�z9)[���7 �G �V��\�sa���k�Y��I�8bDu��Nꍆ
'��:Z.ν׸�1���"q�J)�M�@CXִ��30���|���-��\77��֎Hh�/�j�UMo���8j��7	�yKe���s�͵}R��Tx��)��M)ix�׻Wvȳ�
�����P;�����`�M��|6]p �׭*�m�͛�<�4�6�"��|��LӘ��IR��8ɝ�O1�59Xp��:���F�wj�Npù1?GΛ�S2��@�r��WS���^خ��Qh ���w������dF���fE�-�x6/���)Ԣ�dm0
8D-�l�6��x�k5t��}/����`�Ŵy�`eΤ�/\��LPZ��f@����\Q��r�=b6�BO����]G_rj�Xz�;U�������el�hu�Y��J53ϸKq(P&ޔ0�f7qrYI���N��}��v��8 -�ue�g&�.A�	��� O^�*�8w[�b���9���IFۈ����L���#[���o 3aID�0X_��"l���j���e{��"����/����v�	J^X3�i��%k>睚_99��2����A�<ﰍd��FK^;It���.�:�����i�Iu���������]��)��$�8�|>�B�Da/]�J\DHk�\HިrB>'<&�����R�8O���8��2R 8��,bfu�R}�ᾈ���^I�dS03��I#��X�n�1��Wgϖ�6�?L�/���3�Z�B�i�����O���f���ff_���
qY��!cD騡+x�Zߘ��.�~�O�M����BϿ�t-���YJ\�X��1_U���j;�oƉ��3��!��(���F����L�
���q�{(��~�CX(_{t��Q��K��SJ��۰�4`�
2��k�Q/�P/a�b�ʍ�(��E\n-�V�\��W0^�6��u�5����+��Љ��8���]�D����.�dtC1�
�V"*X����>@��[{�j�f%|��x�EVMT�/ET߀jU���	��6���e���l@��H��r�e?��bƓx��R�y4+o��R���g��E�B��i��aj��vρS ocC�n��0J۴T(i�A��{�@�G�7�{���J0BG=�H;�>]�Ao�L���ȨB�A;K�����F���[��ַ�n�(��v�"��(����>K�'\=����^FE�F�����r�FB*^rIj�P6���L����(=K�oy��pkf��$^�u���U�����Ƃk�Zc�vd�v�ų����#�B����~Os�X��G��RmJ��B^:���\�s���=�8!�b~d]H�z�h/�:,|I鼬P~bM퀫U�X�'��'����JÆ�����?���1?�c��"e1Os;Ng*ʍ�!K�̓F��$�(� �0�̀�T��i� [K|Q׋�Ȅ�Ia�7��^��@IוXD����y��D�AQ�'����<��-w�Q� ��3�S ����Bz��uH���7 �JJ��K����y��.h)k"��c"&��-g������u�b�Fl�d[�Az�]u&`�v�v��~�]���׿�\����1����A����fjA\��� ��i,�5Y��#�	����0N��p��foy���>��q�]&�AC�;X6&Ӵ�c��)�0�G����Vk�$Dh��A~��{���l��mv0z�G]�.��'��m.^:�V��݆�g\9BB��p�/��T5��A6�Q:l���
\׼���4}L�S)���z>�j�K/�\-�N����:YP�|#n NZ�#�ȓSӑ�)�"��6-��.��KE�ᇏU���#�4R�4��J~j��6��WtBM$�|u�IB/C�ѓaz�8�z�mB�3��iۺ@{Y���'�N�e��� l�]3����~�H�y��a�dm+���Dܧְ��j�KG��o��Ѹ7�.d�87i� �`]����f�����f��	�V:����,�vj�0�Ğ����ep�1�W;��dH�$��]��# �4z l��y%k�Tf (�!*�kv5��T�Q����!��=�p�c���!7��!y{�%ZT��=�}��N����M�J8��@���E�g��>�ee�P,���D,n)���8��b>�{6G����~����;��LH��AY�v/���ݙ�'�*+�г>R�_ذ����Ro�ct�b�{�Va��a�h8����E/K�%��{~حs`$;�I�c�n��)<qN �?�ν�!FΡNO˜v.+��(i����IV��tdR�?	#\U>��B�����nM��ů��<�1��� �kl@���BW�K�톱���@��R�L2�W�~�b�u�k�.S<�9~���Bnbd�0avxl�B�%%�T]���C%/��#u�)Ĵ�+�7���k�����@MV@�7��#"��J��Ѝ�Ϗ�2+����������%�R�A1c|���n̻��yR*��^B��d��z�c���r����qp"�x�,�3���$�ʏ�xb���b�0��X=h���T�F$�������i3����s��n����:h�o\DH����Z:��OpK'5��gXë�_R"��#��ﲓ��jy�v��j����6�FA��-�։'�b��ٱ5zc�a�mW�<�[�'�,���S�sSK�e��m���B'�z6F#!�nQ����������"���I Q�>��Pٔ_(m1�
��f(pn�y��8��I�Z�Q���Ĝ݁_W#W���|w��:P�zxtp����[qB	k5���7�҂�%�������c�^�@_��8^����O���ٛS���o����>���!��G��V���_-)��/`C_ڀ�|��i&��PRh$��y<��፳�Y�=�	CH�#�B%Kb�����1�bj�S����"�T��K4y��d�H� �Ҕ�9<��W�� ���We�+�.���˼
�S�{�_�X =쎙OP������bqΕ���GO�V����m���;�tD*��𫽩�����Gޮ}w�'.Dn/�Kշ6�-�p�!��0��m���j���+ B��~��@ t|�w���
�F��GYF�e��|JKzS�����T��R���^ͅI�����R���]X ~y*��?]0l4�P��F��5��|���z3�A�:8[�;JW���Y4��G��ʗJ��$�ċ�%^(�F��%8��#;�k%�T����ɣ��V��xe���d�8��J�5*b�� ��[4o�M��Yj\|���îd)  �� �S��M6�M,�7��8W������(
y���ݯ��$�ttn��Iu��L�h�w͜,f� �z�tᩝ@"��r�?w�D���-`ѫe�E`��k�Ҵ��>%4�ZS,r�N{��hfΧ�����F��X��U�$�N�h�B�U��~���-8S��Y��Y���PZL?̼=cpr}�qc����=�1<����.2���l�_���b#�`�S���L����.�� I��L��|wU�uF3͉֧��fi�ˮ�����k��_G ,����U���Ą�nŐu|>A�5��Šs#<��sغ")��?
'�'��}e2+�12L��I�7E� ">����W�5W�-�d�%�E��5o(�e������B�ۊ���MΠ0W35��Lcģ�6��M�X� �W�P��JN�����1�J
?	CU���)�I��&K�x��!j!�=����=v4��ĭ�I[>	��ټ8Ga9q�̤7���F�K���P�G���-����<�:��_L�z���Z�
��[��b�����/�Og/+
V�i��gFL��\2�7u�js�D�<X����u�� t���>�͊�³"���T���c�~�D$��2h�Xx��(R�����t#Ù����a�]/׽�%����p`J��@ݑ*�BX��T���|SU,�Cb2deu��9"�"�`@���z]�I4��ڴ'�%~j�G� K|���rh���qĪT�b���Bfۄ)�V�� ��տ�p�&5�r|��ֺ���p�d�f�;12Z�>�w�RXj�wb�'MG���{���t�j�m{Q�Z���br�}��8I��HyKvM�Ql��<3�?[M�̇�u<���S��P�ˏ��]��z&��~�Xt��ܝ��!VQ�}�+��	b&��);�q����ᢵ%]� ��)W/ԞaV�F5��$���.�@t�"'�ԟ��>Rp��E~IC�mu#*V���>�ޥ}# �4@��c�`�,F�����$-���q�J��U� ��3���>�#;L�-�M=�P�-{Hz���3;��T^,���l�#����90���}Ii>X^�Mq"��`�'ܬֲ��x(%���h=�"�(gx��n+������!=�(U[C��c�_���	�V�S��)	����^�����Rv<������U�wE*��U	7��@���x2��U��u]a�M�5���`b�?I�/������Ž��d�ҠY�}>�K�B��t��!��AѢqS�gֲH&�uF_��t��ɚ�����.u8���E�%t��nU#����ệ��  ����P�wxG�
A�'c,�o�������&��D���TC���I�/
���������7�T��o���١x��te���T2�X�Ͷ�L��|"����D@n�)�qw�w�][=�_���O�h�zm[��	����v!C���>������4���u��3��	��Q1��-L�e�� �����h��F{T��Wf�M�n�{�lPy�$��$�һ�}�:���t�t���j7c�Z�n	���	z<l�]ZSNl���R=13,34���j
hލ;ԀYZm=ڐ)����������wb��b$��Xj}?�Rc��mX�3�3��l��7w4�Eg�7�Kt����Hߒ�![up��4��á� �(����:�	�^�M�9�y��/����WU1nm���==g�U�!sـ�;��«(6�+@,��OǼ�|��0�c;�[��p.k��S�M$xۤ�3EĠJ}�$!�&�x��pZo���eKPw�L5) �6g�������f*o�%����b��fq
�y7BD���~T�/��%������*��z�9D�*G#K�`e��g���e�9]C�S�����$��"m��mV �pE�f84Y6�),�_�������C�#�|h"��x�r��r!^A˙��|�w�T.|�~!��Q� T&|�S�����hG�)���fn��c,��T�o�CP-�g4hB�*j�n�
��7�f,	_�͕��� �������{��`�D�$��}�}�R��@f%��$�c��=T�8Uģ�����ގ�/k�����Y��/���/3�꒒�%Dd�1�ZW�S�e���h��6z�X�,��E��rU�T����X�j@�o��;/U��hJz��9xOW`6�����x��<VD:,X8��!˱&���S�DO5�Iܜ�[�h�*�9�A�&!
o��2{](X�A _�]g��!�S���n46IE�b�GEΥ�[��H���p�H=�y+	����
3��G����! }y��J�35�jR:��*����V�8Dq
d|+���ä=�Wvr�:~,G�\���l ����V�<�˥�m�-y�,:����Q�S#���A�)�I�� �$�\��0����	l��l36^��LB�|�|I%�ʇ H�P�FP�خ��Bo��h��+��ѳ7�9����6�M�:����$S�'V)i�޷�Q�ꔔp��e�J��s���l�|3L�F�����Hxn^��䪑��jɏ�-����������U	c�xu����?�K� �#`Lg��#��RW��;�c���
�&8�FM���<�-�yH"׶��)$�!��Y���gW�5�Lq�er+5.Q)��T�SN��KuH�]�'�N�蒨�vd*o[�!��	��~t�]=Z�[���U2�&���e�S����&zĩ�@H�c���2e��dWq8��.�7P��X0�`j"��I��rj衫�2�S���vZ8�Kxh߸���h��ڃ��l��mQm�i:�!(QϢ_��3]=���wg��A�����e��z��ɗF�M�(�m)ڡ)a���!���Q����-��7��/�16a5���+�%U|\ȋ7�J��e�_�$#"�<����$�DNf:���1�PH���*�>��S"���5�V��� �A��ཐ!ǜD�__X1����݊�7/�0L>�oӡ8)��Ӵ�ѥR�?�_,y�R�����{�Z�N��s��M��G�����k]��f��[���Nъ���@à������B����gԅH�U5A~�>®w�(*�"��/�[���J�e� Ge�C��)Q�:�ȄC���]�D�F��C�m�l>������t�o�D���u
����R'J$nO*����9�P�G��wϴ�#��<��N`lI6�Z�C���
o�嵫�~]t�͚2&�<5�HC2���'�e�
�� 
�����Au��d�d�,G�A�:��/���<��)��t������KQs��j*�M�l�C݁R*~):�:�w{��T���_������ܣ�X��@0��@�SZ�:�N��U�z�^L���Ӥ�����E�@� �Pn�;�g�����@��D�ѵZz+·�ޜ�`Jێ��!^H��˟�{�a���<�ء��Y_���'��*�pE��Y�D�o/o��=Uh�]T���X���y�!R�����C
u���R���d�IT����}g��y^ۄ��S�ʕ�@d: ߜX%�N+��u<ֽ�l��޽���q�΢?u��*@�jd>8Mj;�Lp�\5�a���Y'!%S�����ΘX�;sd�'��n���^B�v���|;���y��D��Y�"å�����1���] �v>��;P�1%Sټtv��x�f��>�(X�1�R߮�$8 ���ΜSa7���WE;{�a\!�Q�.���-[
�'o�oW��eΆKL��"7";w�R#�����t��me��%*�5�NRd�Ph�X�J�S��:��Xw���b�~Ē񧊁��ӹ���t�Ca�,��kJAg��KRȡ�;oh�`���7��.-
�k�`i�f0;�A��,��O$u���*)=����<�!�[�8�k�t[�����g�T���%��6¨���T|C���ff�؃!<�b��������h��I����k42ؚ;+�0���rM�џE+�5~G�|	`���")i!z� ��]�c#���0�6�rĽ����u�ON�ʺpr���shv�/�+=�s�f}��:�!t
H�I����:(#�
VS�����P�Ư���M��� �����QF5������>�Ǜ���,��J��U�������fSQlP���k�=Q	Rk�y��ר�D����� �8sK�9@�X���ot8��j�����]@���	Y"gOv�KdvB>�\ϝN�#1Op�� �0����O����u��͡~T$E�XDj����Ya�PYˮ�^��e���G�|bX4����˶&������	��I��*)��\��Y��(Os�e$�h=<���25h ��3L����˫����A�փ��KZ����r�2���#ţ+R&EY�v���Hy叿�&��2)Bd�68xc}̯<(�����)�5�(S�1ˆ�#�+z̳�h�f6�ӛ�D@2�lז.|�l��!JS�������ZPY��<���4�۠ϑW�FY c�.�'�#�@u��[ܛ!��"nX<���O�=���?�N�+y�S����l��m)p)� X��k~#SX��[FY���9��5KE�w��7�F���otIg���$�IEaeܻ��ٵ�'0�tb9޸�#�c�gǄ�v/�}Qƀ��(A��3T;CQ�fqs�:�V�oa�՗��G(y�+Ƭ�I|ɩ>	*(��߰iњ���D�Q>�����N�3[���fj*k]��m^���p+� �i�����U��k����\ݪ�j%�'"!�ַ4 �b�>?@Љ�k�l��_6�z�Շ*�i,y�}�̔/)������w�4�N���&��و�=v��$H�	a�m���2k��*�6��N1����$�="�}>����y�C�S4~
ax5d���_(�6�#J�-����ַ�|FDN�:���ߪ��65����e���f"�А�Q}��b(��i+�l��l���q����r�� ������E�N�sr��&�!�m6kJ��4��Uq��P1�p�wY�˫Ր1�)0(�쌉E�s6��a�����0Y2O2�loKd�A3A�����3c������c���%��Tۋ��i�M+��,o��t�9�x�{zo�-��d��þȲ�ǎ\6=,��*PW���\r�p=pF�
*7Y�r�Px����c~.A�;�CI��uQ�H�N�ȁ4:&��v������tL�]t2���������Ӯ��r��������;��#��,��-����:�����|Y�,dER��a�,���D�H.��r�X�K�EKG���9,��r����y֦���q��>���I�j��9aE�F��`��
H��a;L:��A}��|a F���ɐ.@��A�d���7�h#��lT���"�����^�������G��F8n?@�wFyt{W /�����W�l�R)�y��N��t�iTo��`|$��OZ}N�R�k ����	��j����SܕK�,�&{��4&T=�Wq��il��6P����F��K! �Ot�?g +��kY�i�H�_�wqk. Sz������+�)�u��[�PET9>��!v�r���?a�d::x�t�9<eRd�	�~�_EXےP�w8�ߵ�
_�]J�߲�j����8r�v���{)��?�<LVG4~9�n�Ơ4RL�b�x�w��Nź�pV�G�;�?ې,��j��<6$d@pnd�&Is�~\!�0i�>��<���4���Ȗ �1FHmQq'�P�1���n��O4|�x���h�_Tsڕ$��b��@�yL̘�ƅ���#e�4=�4��pix#>����|��0OT*�sDΟ�a��5�6Ŋx�V(ԈL!����^�B�f�ؐ�.W�)�r<�|o{��H:6�����@��*�ʒ�>O���G���p�T�A���%��_�Q�J�&�m%gE�e��tw��#��$�v���8�wy)f,p�p�D��D�afu�k����[t���a;�ʆ�I�&C��Ԭ�ݾ��B���}C����V��t��Jc�M�Sl>����,��.PF5�o�{%Ļ&ճ��yS��^l1�ݳ�9��Ǜц��4Xږ��@�>��cM|�#h�|,V��β5�"i��)L3��:C�:�9뷀zb@ɧ��"lƞ4���mQ��@�mY�@E�`��ߚ��:	�c_Ǐ��Rޒ�'@h��#0�_������G.C�G��ɕ ����?�,��\ͱP�o�dwaV�OV8��-g���Yߪ�W(6�\����cf@+�`��:Z�&/��k_I+yC$��1�RF����ӘaT���+�Z�`��r�F���9�L9�`VF~S�;]�rh�D�}�6_jfs!'(û�, ]�Ib�~z�6�یV��O���S^�q��`�ˆ2�r��AJ� ��޵DL#B,����5eD{W�ר���Fޫ+\�����쬜�d�`zy�����;ͅ�i�e�� �1Lk�'O���$U�Yh�O`�D_��J��/��=I��Έ��;5�ǳ#j��`��D8jN�9��gf*�)��{`��]���6c��;y5>�9��K���W����M^ �&M{�܎Ȅ��1��0LL��s?᪶Es��-���ﰥ�W-'��j��=�Ӱ���F�g�3�/��n�#��\�D��5#b�����!L0Y��KF���a>��N��!C*ngN��Yi^�$���WH1��@�]�ƚ0���{xR~��ʺ�!�M��Sx_ت?#����v@Ԥ��U�-? 5GFt&�9�I~���#�H������jt�]��g�/�����h͠�=�LJ�Z����n�/8%���7�,>�q̞��'<���/b7ډ�'Ch�N����dԇ�>��gd]{�N(�+���GӸ�^9�����a���&~���#.9��>yY+�v�Y'Ō��R8��7\�N��\�A�H�N�u�k�RZQ�5��d���)Υ�^]h�[��S*�)M�G����U����h���p?��E$Zw�z�1��;�>��x8(�4��yI߼��A�O��$"Y M��N�<}�`�?]��b�ѦG�>��2�w��X����г��d���DG1U��^TZt�9d`u�$*�B#PF01aEF�s%�����.b�X/΁�Z)$D:�S�|�FM��/�l	�d؇HE����v5b�����JD�����e��-m{�s9 *���B��]��@X��%*q�����0����V�Y`��f6!��d�gr�̻�J�@�*(��H5t��Z�7���������f�ė�	4M�.��:>u<�I�h!��_�I@f�*Սܝ��DC�E�S�৙�	�zߡќ-i.�Y$qc��C��9^o�J��˞�0WHVD�p� ��r�^aT��L�P��k���@�rM2����zw�3�M3�wւ�s&0���1��JEy�A���.Yʂ����;0�N�|�
��<J��l�z}���!X#�d� �tb8A�	}��BY�!���D���b@���I��zPR�$��[��.�<���^��
�nJ
[tHϭ�N�����?�����O�Y����d�����Ig��i����b�Muc��m�3�Z�ez7�EG�z"ra�h�� �X�~��B	C&G����8n&���d��[�pŝ� �1���x �~ī��X�]���O�=}a�1��
~Ɂ�C�����6�Q~J�徽��&��LN��}O�^�Բ�l���r�iu��R�tsX	l[<Fɳ�/ڀ�u��2N$b-�|d�)/���Z�4Tb���3 Ő}!(zv���`� T�h�4�]?�yHjRX�v�Cy���u"^S;"x9�
0"�PjQb���Uѯ�ָE\��S�<�Q�$V����4Oa&&�6�,Cn'�X��@�,�T�3��Ӟ@z5�O|U%o[7�'�*{ꂹ
�x�Ë)���%as��|g[d���pE���U{|V��E  ��V�O��x�:���3�n����!�#B��a'"��f�,��f�M��Ұ��%1�0�*��0O���=	�i}����i���Zڑxp�Ř�zqY�?�擄s9|�P5�
%��L0�.4>�5�����	+����žzڎ���g�� ��73*'л����tO������߄�^���w/	��#�j [ŎX<��C���*��\__��B��П��BX�����wE�b�
��x���C��)��3�%�QV�����J�|� ��q���fi�Z��c�gt1�c�,]� 2�%Q }�p��n��rT��-f;Qv��2�D3�&�5� �1���)�@;RKwgU�>���\��S�D�u��b�p;U�*C�tc5X؏-e"�]u9���!�@I �r�|��0�����Y��G�
]-�d��ff�呷�
��I^9�����#��(ܩ\�ѶA�U>���̠���T6�0A���R���D���X����R��`��sZ�d�H�!h�lJ��������Z����&�~�H��"�r�8�|@���ӎ����:,�,p�<��O=�Vl%�h�J�sG�nR6��(&�M��|�������oI��Hb
>5�&���������uoC�G+��=OW;��GTz\�G�����z�*rr>�k!�F�*�X�?,���a�RƢo��6����,���l�����9�=��w�lb��	%X��,�tڲ���.��x�
f˷���i!�vԐ��uCԘʞ0ͭ�4_ɡ�c~��{�a�:�|����4zˡ��'Cp@�x��G�����n�{��F��Ζ�Fr�.�r���,�nT?��JѦ������t��]s��!�eۻ�.�N�I�\�F��-p�*{���,?z����B(������1�������o������ku��&)㌠P�a�&����q�g噸Ϙ�2X��gB3��;��P�H�Y߇E�M��,����k��n�(nkS�5Z��P��u�շ�O���+���&�^+XPO{ng펥�i�4��"�����B��ꢤ�qD[5t��V������|��o�..W� �Ͼ2k{��z7�/�->y�S��&���-|�Wb�*M{ֆ�_��0-N����'��)�����|i���P�s����1MBh��� $�?����R�&ەv��I�.����@L�x���Rز�V���iԜya�N�Ap���d���e$��������q�/��;D��g"����φx��|2'��E�^d-E�����3e�������t0L=�k��@~m���,�o���1���De-Z��&�����vqpf�B��"�Y -��UH��>�S	~�J���C�n�9��/��s�й+�c�?���$}pq����|W��s[Ť�!mu��������y�t���.�g�_V��-"d�t��J4�[m0
i�}7���(%@��jz?2�����c�D���n�D�]ON�������E���u�l�����,_��Hsś��ߏ����[qQ�c���uU��}x�Jj�e��_����{+[N���?'W;��+�Zʹ	\=�eaRm��E�a���dw���ʢ�*lzr�v�0�Y�!�.�-�����:r�}0�`[�h
�>��KӸ,v&���y]b��&�6�j��D�W]��?�W~�,��8^�^ȉ�V5XH�c&#�w��ѻ�i��U��;UB��z�4�X�v��lY�=Y"��HlE-�_��K�kp�1�]��:��:�h�
-�b�X4j�����s��
��B�Y�#���B�m�'�˱�6��5S?��! �n�����Ue)T,���	�5��rTN�i�g*[~�K�Q��������㯒�W���W~f^���Ѥ#������F�zԤ �QZ��EQo��X"��&�5?�jF��n��.YF��pŚs�#�܏�?^�iM:�c`mI�f|���˜��������a���Y����d@>�Н�:�Ώb���v�}H�C��_�`M������ͭ�G}����l˙�"��/o�K�϶,sta;p˴k9B	���P�˦����[D�QC�%J�'�Es�G�6"]"���
��� �J@���hN�c������B8��κ����{�lޅ�B}��$n�'�JS��a\�I��9�3�#8�E�&"2�yMװ��q��j�9�x$�Đ�[kbw�h��D�7����FXY�'�j�F�i$w���� 4ѝw��Yb�'��U�1ᶿ�H��� ������&e���Ar�ʒz�Q5��xj-z�)���
�����e��h`9��6�4zzF�N�&zyϝw��w�6py��HC877��;�ݞ]�]�k�����Q�R!��2�1FU���-=@���)��(���<G6Q�
�7{''(�*��CI_�0夲���>�j��R7(�l���g_j
$�*�ce�N�e/�S�����H?��-��ڥ�f"�u}<d<]�1����+.�~���/����y�|�c+�� ��i����]v���)���_bv��uǤ�s�UD17;8�zkB*�Nd�@͈��f���ɺ��6�tRO�<�s��9�HݖBaU	��x��7i/��+T8r(�L,#�Z�x`�j"tߏP�@9���b�����Y�6���6;m���{}�T�#�Յ��pb�o��Ш���ꪖSՃ=H����(E�L�bg���,�y��&O>d��k4y�(*Si��F[�e_���x�ޮ�:��7�+�I�)����|�H��j;�y:Z�M��i��u$,��|!�%�� 7SqT�C����:��3�@;$���͝|Ci����;�K m�j��������6m�<��}2�C"�`�1G�Q�`͖�2�M�a#e.���#�T&b�X�\��I3�ɏ��:�m8�J;�$�~G���\���)��k���Vȷ����eY������T�A��L��u������f����>�b�˭�??�P��.�1��~~���*V=8>� �E�$�꜎B���h:A�n��M�NKc��$��l���TEQGr"wX�ք�,��Npf�Ҵ���k�"��)��{s���S\���`@/�Xqٰr��F�8u��$�:�< �������ڈ�B�MA��	3$p���Xg�~���J;�T��͋=?�b]�c�����s�V'zj���P7
��g�oȆa_|s8����d����<�"r��/����K�u����"K�h���T��cH�|�v�uȈRY������@+*F�z"�)O�z��?�Y��.դ?���'��^f��r�Y�����.&"�*�YS�{`W��H�t���m��f<�Z*/���*�R�F��o ;�B�
�1Q�~|�%ek_��~&|���o!E\`XQՓX��	'G�cV��� ��"xBu�ߨ�Fqs1�N(����<�%�[���N�L���n�)��hbm�T��7w��~bWlR��k�	����#�i�r��)6������{��:�7���y=����qˡ�aЪ�۸�@�Wk4`�V��у^Z�yg��e �:�֧E��΅�w���I]��=��-)X�-31�I0� �x�	o^T��"����d�����h�ef�n�AV����~$�/g�ٞ�����p[�=��<G���s��3�i��q�Y��;"^� �^�5�uca�b$-�� ��O:����R{w�^ ����r�3BG�O�zF����
o[��j5�nD�qPe��%��0�Z���
���7w�]͆8���F��<���=�U/9{L;A/CaV�J�ټ�ՄĲ"��A�>V�mH�<M+)_����R�Z�a��d��F_m'u��q��3w�ގ̖77�i_�I92C�=5�.�*���t)/� �T��ﻉ��x{ؖU���pa�::�p�Cd���d�{ӊs���4
�ͪ2�pOl l-���/�RKQX��h�ꗎR��H];FD��	Tר��>�MJ�W�G��T"Be��.j��eRA3��=�)0<��4��p��|t}����Y��9>:M%�[��]��02�d-� U����bk� �����ev�����M7?�ϣw4�j������y`��I��GRJ���qi���A����}\�/L����Ӑ<�=<��X��)5B?�=�/j-Ѱ*Nm��qg�{bHֵ��=����:���Lv�X�G����<�F"}��D̛�v�h�BOS�5�~�%@^ �V�s�R����F�'��2d!I"/$d�i�0;lR���Llݑ��9r]R?��5�D]+�$�������z�$FOX��25�}>��O%�MY�"L�cw�r]�F@yF �=�� ⮩9��B��nx �h�Y6e�R������?��S���T�='v�c���+TiQD�煺��.���noa��q�}��l�wp[*��q,��/
�oO"�(P�-`C�u�sy
oN;�}��'�Ւ����y8|�|�?��O�;oq�_�Cxm�߭�x�82F[�Ħ�hB=е�\W}4(��%t��Ԗ�Г�(���� MĎ�%O~��2�#�����4�k&�¿5x���& -���))���ء�f��$y)Qk���G��X�L&��J&�B�N#��F������8��Oi=��~����~�: �������Ģ���R
�ݞ"���'��	�����;��e46��E8�k�Gl�p�����T���pR�czZ���Z�!=�aof��EOT��+�h�i/3Ғ>����n� ��9�/��š�WW��8#�+����	����Te ��q~噯�vB�� ��P˅�R�F�?Jx)���Q[:�H�7���G�)���@���u���͎�{7�G��7ɨ	��q3sj.mؑG^�θ,�Φ�%Ď��$gU��$�[��=���F�wY{b�e��2%��v�ޘ���cf8��\�J�ۢ�eZy7��}�p,n�oݶ1y�@\F{Cs݁�?�@�=m95[���#8��S;'��:�K�`va-��g��&qv����A��e\���*
�״Y�+"��L����
�=��3ѫ�o�{�s�*hr����C��|uxdx�Q�غ2��$I�u��Ш�a�=$}��CI�'aՏ;o��ι�V����WB���C_:�-F�3�R�T�S�t�g"��sS���8��O�W����E�aM�?�$D~]��c�| ����i����:*E~�J�������_^�}z	7w��&��7��`[�V�B�T����+��
�*���\}^�alW�#�%��"a[�w���Q(7p҇�E>��6�+�'�N�H��^�OW&ܙ2����zפ�;��ƣ���nk>Ar�'A�0�|AS���۳��F]"CKl\�ǆ&�'吡
�����U,kK�� {�g��%�ԹO�K��g�f�1�`]I7�t ��� ~���m`8L��u�LR���lѱ�x
~�L��`#�*Ug���(��z�v_�b��cDr����jLV����V�T�w���;���x����蓳5%��18�)
��8��In�7'>�|6�?g3���n�r�jI�-*�(A��-LMiǲJ
П�@s��ҫv��~?���t�A�q��9���Ųi*<��w��Y��Gu&>��|�D�Ӆ{�1:�a������B_P�.{��	���X����f���h���V�E�Q}��R٧��Ӣ4�x�k���A��;D	�j����,�.�Ӝ7�e���s�^��/C���Lw�ӡ�4���k8:!����yS�ZkD�����6M���ĭ���!>�b��*�̈P��=�c%+�G%9�����Zf=�����������.;�5�:6ٶ�1"�=�b��]s9,�r�e_�ٿ
��Ѯ�D�J �6�v���?�� �/��3��Sa�=�X�A���Z�{��|�+�V[\�囅L����ir<�ud�@���k���
N��Iq��a�V&��YI�ЊD�v��ǳ�0۲1�g��2U�d� �\C)���枩��qSƙ֊����Ũ��1R�0�wԩ�fӃy��@��Ṡ��e��t����v�Tэ�z@�2�y74h�7��N�n�I��z�ݐ3��T��¹k��a���p�f�ɘF�zh`}����0�����
@I�YkR9R�2��?bH�1UR�ݾ��8�'�	?��3c�*�����[���c���d �ɡ��%ɠ�O��/Q�*&��ğ���\�fNBϐ���2���` s�c �Up�Ł�B�M�uL%��#��=b�"F��v[���Y��I�Jx��¸�X���P'���du����"(|�`��m$��lv�>��f%sI��Z;��8e:�#�S�i2�]���$�:ڄ�ƶ�4ٶ�p�bjz�OQ��qݐ�U�;�T���(���A�6y���lm�~��P6����ҿ�_Fa���;����(+Wt`*G�g�D�6�͓�y�7��7��1�ݏnDg�S�_��5X�̽/d^���v�eM�v�sbv��&�	*�R�@ض��Y��U_r�c���(TIR��>}��5ӑP��ӛ�X��
�8����&��q7�B�t��G��O�N�6�^R�i̪B�D��R9$k�o�����+(�S��o/��L�H�R1hpX@S���1���`����]����"��lb��.�T'�,Ͻ�T?��f����~�=�T��ռ�A�)��̇�zE������wk�!��r�\�kB�,�<_�����`��xJ��W�K��+�0~�}��#V�(7^�X�h�f���_���j�?�vaM
.�b%����,�+�e�������mx"���f�� �/�$أHH���w��?W���CD*��yU�m?�`�������=�,�����鞰|����Q4�'�BАC�g�-�O9�+�[0��m���N̡4(2w��)`Aɪ:Y��2^�KO#�~vJ��Ej<u����}An��!S�uW�&*�zA>�m�l�(�.�w��&6IO��#�pž�����"��>yH���4#�v#���e�,P�||���\����8��i%��ǂ_\��	F���ւ(B�����X�9l�fߠ�x��?����v�v҇�9�7����n�X�k�����MZ���D���|��BPDd �\G��/쭽�Ú"�܈�D�]d6MB7��VhY#�q�`�r�~80S��b\�h I�Z|��!�Ma!��Inq�WȏL��Dx`X$M�\հ+<*.ae��~�'���� �ݚ�K���KդY�ӳ��y������Ytx�B��3?	rg��Z�?\�WU��]D��l*B� �8�!�yg�����W��ON���Z��u>z�քk�w-Iʋ-�?�ϡ�(����h�i�_j�^�t;"��C���B%F�;?�) ��R����'�&��̖,�� Qp�O	�߁qF�
5C�ֺ���6�l���'Wk��t��K]1���{7�e ��;��/_�n�E FV�h�b-n�?�0�/��V��9 WԹ��0��
A�,�C�������z�����F6h-qy�$8h/f$W��`1���Vw�<Ht��;vdq&�=O�1��X�[�~�@��;��I�_��R��(��������{���~پ�>9�Mъ��稝�odîE�2,�wP�]� "��E�s�&i�:(;~x į�&�5"L����o`�B�P�ؐ:E����y�j�c����`�@�h���X��Rep��C���sa�N�_%����
�6�)�U�oO�궟���|8Ӛ��S�KGy�p���sZ,�9@*��h7�F�w�^N�8{��!
��p���Ur�����)���1u/�G�|�f;*�ѩ7�]v)H*��%���d_5z!�M@�Jq�팫�fuȞ;�+ ����1CQ�R��1�<ޒ�,����Z�A�\�*uvˁ�\C�88�Ơ��O�>�~k>w=����q�V+��c}i0''�`�*1ߺ�_/�>Y=�A�Ǩo���z� ��_�G�����v�d��is�����;��L{<#	�1���M���qH����C�U�aܱ{�h)��� ��eP�6F�!���\0#߭r��/D6U;6�C�g�]�)w�)jg�
��	'߿�D������b�*Җ����m ��8�f��_�E�Y� �!ƭH���He��zmG0��,J�Y�dUX�9?%��.��v	3�+<��G��d�v��X�(�R����F�/w{�}6]G��U�ŏ�m���.{��3�=5���lc2#+��p^^,�g_u>.��f�1M	�i�s�{.[MSr�H")�V�p�OJ��m��
�g�}ã�l�bNW�q�AI(���9���nX�щ�t�d���d���%��Hc*�w�Zɮ5^�&��۫�UG�Nc�l<��
+������ֈ���<9��L<If�G4�=ۜ�6���-Jl��bO�sA	�E���\k��T�,�o�UR�ٴ7f�r
�D���eт2/��b�ׇ�����k;ovv����s�.*J_���s��%J�&� vM�X������l�'ކ���=��zYA:iw`�%���3O�O���)��J��-�5�g��}� �`x�Q�P'��]�4f،J-j�qy���T��e��S�~Z � ؾt�g�T�[�q#
6t��㧨6o��v�0W������k�U�O��C���>eй����J �M����6���(ٽ�W6E���bwB�Q��B�n�V�q;�BP�R/7��9����Z���CX[��ק�Qб�/)1� v�JU݃8�=�8K��iG�_~F��QF�A�r �'S��05W�T�XOR�X�c�-���.K�v`a�'hG�_�G't}J`w���{�=jlv�2å�Ϭn Ő(�M�S��	m��F?<V��H<K��5E"�`�C	�=5�G�S+9-.4�.+Â�]�.%?��*ɵkx H�ƫ��Mf�:�������lp��M���	gK3X6nu����T�� �7�,����E
0m-�u�S���@��0%���n�%�����8S�@!�����ՠ\�����ʬ�u�-G�¶n	�Z����Z<^��P��A �*��^7��}M�����]ȅ�3N�*���fj�Y-m�#��9��%N��1:�ek��`��/Z��I�8��=Ҹa�Vrz�<ր鞞N�b��C<9����KT�����W}R������(n_ܲ��
i[H�滞���oX�<4s��'��E* |3�� X�+�u~�a!����8>ؖT0�*��r�� ɴE~d|�^�1��"��c�D�m�t��������Q�b��|�$���X�zS-��I�02�Iqa)~�32��ST�:��)��ϒ��9�y4��GoF��-qR��wx��78���)J���n	�-G���.O� [(Wa!򫊘 �����!�$ҙ�D�FE�m6��;��@P74ΔaG!�_M����*�薤�2w-�
��z�LE��[$
��}J�co�X��3z��Q�;t�j%��|2��R��� ��z+�v�~B��p��3G���mmfɴ��O=5\�(�]��`�H�����?ێl�Xޯ.<����%/�7iY,�bۥF}��7�x��'���?�Ѹ��҆��<�v��c?4F�Q�4@'����
D��*yH�y�4�`�O^��Q|Ǟ�;BJUS�gM�!}A �t ���6GM�٨���
چ��J%���`2��O��]�È@�=c\d�d�|
p�!d�.k�:�ɑ�_}�|%Z&��cA�m9�g(�3�ɠ��P!��7������z�}�	�7x��6�`Go RX�KJ
�F�U8!/���:�&=���ϯ"h���`�E�Y;�󓟋h3k��+T+�❜�!lU�x���\���4�4�*-i3�W�R,x�k]�i���������.�±�P'�=O��{/y��t�O�w�%�Hd��B_��}U�؀�F5٠��KF7�k4D��E��;	zĵ�JS�V�[K������ҔX�hq٣��#�m���B�Jp��_��ߍ�2"!-�~ ������F��ǧF�s���w����Y(�˾��@��.OĜ��".[ͳh+4Σ��g���F����E�>��5���ߓ�E�,�� ڑS���K��K�9��C�����L*x��^T0�}�]ָ2�wQO1^��mu�	�z{�^_{����	'�M˶?!�����P�ʔ��U�:$NbW8��\����¡�5"�[��Hc�З�~���R75��ӛ���*!�0UgW9cå}L�˺d�j��:���%"B]���F	�@���uf�/?���H&��@��QF�@?�\�Ԙ�w=��1��z����ݍkun@Ƌ]�bCx(\z���ӏ��@�u_!�ћ���!�h�%����鉢�柹"��z����1�nBPͺ�j�5��2~}
&<������f���
�*gn���yא��)g̓�[Q�X�3��G_0�h�د"�X�)���H*�)�T���5���Q��݇@]��b�O���_����r��U'N�WZdl�v�_Z�mA�Z=H4��
h	y�yj)��&�*��n�[>����{rWX���>��p�F�}�'J�z#�(��d��(���ʥ�n�2C�M��8ϗ3H9K"�8��A1/V��=Ր��r�E�>b˼�S�c2@�I�3�{F���h���-\��h��f��ѓ�d%���\}'����$A���ʸ���_?<D�������]�ҍyxB��ʏ���s>��Nuw\3�0k�&��Pr��A2^g$�����ņ$�^Jᤀ�2~x��6�ދ�k��	ɛ� �?t���f�ٯ��K^��d����*O�O�I��2�+V��'���+���;U����a%	I��ElqR�eUP�P����^�5j������"��XG�C�3\Gpuv�_i��T���䥄��{�r�$^�'1$��R�ȫH���Ɗ�e��1��r� y�NS(��\co?QgR���F����+)A�gYa�5	EL5���Ձ�J�a�T<O
U��O.���uV��Lu�iW�3=ھ#KnY�Է1�D��f�CF�/�M��mS����r; �K^J�2�1��FY�o	���>�j��X*L�Uz�o5þh���l��<\����@һ}��X��̈�' �|�?���E4�Ɩ��l6k^�`����)��(K�_�4g�h{w��3t
����jKC�w8��5�<>��:�j�ƀ���36��P�C=1/��6�v��2,t�j"��w�Xx:ԯ'���s/0M�7��_!��6��o����p��#���8)*Ts+��k,����R�Xy����h�bz.�.[�[�C�+`z~J�:z#�����Ł~��ϩWb"A�+a���i�Gar����bk�x��\؍�P�x}�g��>�c��R�X�Q.���r��|ya ['�# e(����؇q�y���{�XcV���B.���4G(lg|��X��Ŭ��%0څs�2�����u���H���o6T7o�nr=�u|�Ǳ�֕����"5�W� ��4���.��F�u�'
t�Y0����U�b2��)�1��O��jC��ר\�%���>�+Cskv�-X'X��B�_�H���1�݋����Xy����a���m�#qz��(E�5d�*ҴO#���@�O�v�gvJ�����.kEZ
�N��6,�E���E���:��S^
�gd���h�;� ;��z�Cn�Վ���]8w�	Nv^$����2h��c�ىO�D���0���Iƴ�;>`Qn���Pek����(��g�~wH����-�|h�2�=]���$7�W!�K��E�3+a�Ɠf>�s�G-��BQ��f�B�L#�P4�f���� J��\�㑜�<ǣ�k�T>�����qɺ��)����)�x���ڢ��(?I���*�wv����̥�@�a���?�U~�P�]���Ben�~����Ό��9U;�i���+�uF�G�w�Ѹ>�,�~�8ϙ֨�K�!�E�i�gNˌv��ה/U�rNyک�n48�-?T��,Gb��Xvǵ��Ϡ("�b�JM_��@\�����3$j ���J~�O�� ����BuFOJ��zIh���c��Ͳ'�N�S�œ�j)B��ZO�u�1Ltqþo��[��}� �Ԗ�ؙ�=�R��C�4��}�x�t���@�j��WS��΍s!�J�S"�V����Tu�Gث�i��F��&����0���^����{���H�B�BV��H[صh�m����3��f?��.���Q�wh����<}ޘ=M /Sɖiq�ʵK&&˞������6�����?����Ӿ���nA(7����_?G��8�9e�f@j/�t0�8:_~x�h-7�������\4���D��;nW����{�'�ک� H[s��Q���cA~�k�t�	��9��D
�2`.+���܇#���%#<�-H��VZR]�du���ID��s�߶�w��b�v
���@�.��y?��$I<MKHu-9��ѳD�_���f�*�����&
1�m��+�r-Rf�`�E{j��\��]Q��y�Xކ�����'v���[+w*�d�T�IIBb�W���=�|o�PR~����%	ʑ=Uv��kZ ���lI�*�k�A8>�i��b�?s�OBׁ��Dt���l�\`[:P�Y�������v��El�T��,���C ;�G
u�k5q�/VzF�ƍ	h�c=�fF�9ۇ�A_ �So�]L���Hj7�zg��g��l� W�a}^^W��s1����=�Y��j�R�9Y�Rr�=^��=J]K��,��*6nG���_�n�zHj������v;Ej�d�"�\��Kr��ΐ�Êk�R�]�P��tSf�y�AԚRP��Y��4��3�=Q�Q���%��(̊oV%_�	)���<L��;("�?�Qzx��2�X�l�S�1�:$�؅D�q�fG�Mu5o�-@�K����׀-�?<�$t�r���䶳��ɧ�]�X�Cp�v�Y/��Nܠ&�R�mw�m׮ҟ��N�=k����4�1�}�����x��˗�0:	�Hb�5����%;�f�/[T;(�6!J8"a�J��?ŃF�.E�'X
T��p��`T�&�N�˾?�Q;cC��pO�>�X7�	E}�
Y	+�f��#�'�	*��e����<6U��n����<iZ�s��C��qF�!������s���2� BC1�p��e�5��>�����m��H�K*�A�p��?���w���)�W��)OiX�		j�6����^��;���gE��˞NT���A�PM��XQ��Cm����&9)�ɰZ<WBhUg��7�)EJ��:a�6kz`_T�b�4�AS~�d�Nz�ك�k�C���7��P��F��J��g�	D�Ed�K����Z1)޾���Ti�D熔5paҩ������� �6f������zp~}�[YzP���4Ю�U��m&�|�-��Tx+����.�>_/U���1,�@Ѹ�f�zЃ��rsr�r��~g)bx���c,���H��M��7��m���Ku�i�}���W��S*����E��>W3ת���_�c2u/�"�k�K� A��B�a֡��j����*Rb��QP�b7*iL�2i��Ԙ��iE��x@ŁIͨ-�3y|([R�~΁UI+n��43O��>��4C+dV-��Ь�k9?ށ�/{�;խ/��p���.�cR'�8�,k1��\f���Ӻ�t�N�.���gJ>2�\uK��:�÷��E#�O�k�#��9�Q�@X�o���S��
cs!S�$�a���uRɔ��������IU�b!� >s'>��y����V�=�Ry��"�g
-A0�����;�v��y,]T[s�.?�}���'�N�8q1����Gh�X����'�\k�=�s��X�9����u�r�k�[��sX^�%�oĂ
�^��(��N�q�u��.�q��ǁd����6�����p ��7jo�&�	4_�<�$�t
iHK���p]����ӊILu8ae�$cexHi�6s�F[�7i�!�j�Cн�-V� �"�Y�j0!�����ex�'-����u���P�I�A\}|�a>��J����y.������o�\ܱMo�O�g���5��ʛ�[�˩�-�b}~�n��&���u�=�o|g��������y�m�ն�W05��re��t�U/�Qj�F�/'��iM��I�&-vn���4��Wd~>8��d�w�(���6L�d�׳p�fz��@T�l#[�1��ӻ�����^��P�|W�yLm-����[
6!�Z��-�@���]��y��	,�An���٪c�o�Yш���X�}Vy��+=�|=�Yw$u&�\5�� �T>��Wd�;����~�گ���}�o
��7�[�I7�'��*! ~�� ��!7/U�xL�⇰�1p���d6�a�R���/=���!	�ԕ0i��e�Ԍ��.�2T��J4��@k��C��CMb�M�٤j�T�?4e�����Ga�f���_82�J���ߧ��p�����f�,�-��&�L.	Sf}�Y�Эp�����tWl4�s�lpM)̽��$O�0�T��$������Tʌ���G�Vz�^!O3>Te=e��|#���S��:d��x����s�ִ��W!0���C��c��i<�^k蘊=��ߦ�Ž�!����X�)��%�h2'J�soL����n�9I|%�.咳�&;,w%u�=e7�ͩ�����1�6������P� x�mࠋ�0�d���xB�ǜ�m���=m�
�� 䋫ڷe�;�Ly���+�JUkQм6��!,Y1[�=?6罯�C�w2#h>��~#�#�/`��t]'z6sZ��[�����Sw�!X'��=��Br�(b�sNTx��ݚ�2��]��狗�
Pٔ������d���zn����éJ����y�G�kF��IM�֎���4�#�:�-�x�m��+ә\�;-������K����A�����o����*���	�E�16�Ч��P=�a'�U�����g��}��n���09�SL K�~��͵���1�k�nGT��1Z�3v�H�t�2Tz+�C����#彴�Ҏ>�}v�Da�2���ͻ�,։`��s�Q�p��7f8���ۅ�.��Q�l���L�`�k��d��xo`�NS�K�X��f,�kdwPz[�!��M�44l;c��٢�aQ�%pM<��S�����@^>�����k��g���KDҮ�[؁߻�ORM
���O0-��\�u}
��]R�E4q�n���7,�ߌ�]��(:i��g÷�	#B�{���@�PEγ�Mt�e�*N�3�@ڣUE�'6z�aQ'լ�������?[`pdA�c�����G�n�ZfKS�J���/d���b��#�[�:�y	3��f��B�W7v���:���fnW�Me�-�����`�S�Hgy�L��0;�j.�1�rFa���;C<�J�6�]��,x�w@:�]�$a�b�K`�/�-��ڨ*��5 }�,ߵȗ3[5�H/x;K|b6�&9�fx�@-E;�yYE�1fk�y׹܎��^UROE"Ӵ�nP������1�9��ۛ����5)���V"��D�Ÿ/~� ʱ?h�ѣsE�4��i76�.�ϖzK+H��1C��WEwP����;f,��}��U�@nI�n��Hdۍ�d�� ��b��F�U�rf"jl	ޞ�|��}A}v���3�}��8��A�Z}���It�ا|��mfj��`R��5�Ld2����\R�Ჵߩ^j�+���g��d �K�%�*�䚠L%�y�+kɁ�b���Џ_��* Nw���7������֒4  �dN/X�'t�.�2���m�`�C\��5�
Ӳ��7G��K�ai�sTΟ�Jqh�8M)�X�9n�U���B�t���ұ�a�R8��}G���F��~sU�K}�|�N�ռ�C3=��ߛ�&����b�=���q~0����<���dz�qL�̮�.���I�v(��g�Hĳҏ%�e�k���1q�E$}���6�+Yކ��_M	;��Bz\�c�<Ug��z�H-r��oS�/#KǤ�Ej���*��?%�����`���*�}b��Q�/��}��?\���$��bF��׮8��"x�T2y[��9��NΗ�#�ӆ��!K�N[?�@}qzј-�m>��3{!��7�cbfm`U�U�����gl�K�����"t3� (�/HFIr�3[�!)a�r�+||U@��-��4�#^2�����[0/�Cu-~�ڻ��E{��ވQ�ȗVA+Á沑��j b���f]�U����r��Ip��/�MW������Q�XD�A���r{@�X�8�t3���+�̲gGcB�-�K��Eh�X���Ƶ�C�=
˦E	�����qVK���4������O�p@����x�Y䪮
�?+%�37)ƫ0�� �E���=���׼��Z�{}�tr��MA��c.~�Ҙ2���	5�;�!�*Q��B�R�=R�ޢ���t���L���	����Rƃ�UL�o��);��>�.�����?+���e\( �h�)�($��w$�5���]��-o8�쫾aF37ýc�$�_� U(��V��U��%1����v��M���1�>�A0I�䨄)����vɟ	#�����C����ԥ)\~-�f�3�1�$�c��X��W ��i��;yco�5|�
�*��b[�;I�m��hA(�g�e	�T��,S�A�S�F9����B�U���[\|�7٣���*����k���D��̒M����D�/p�=6R4�'��t�����
FQ����@Y�;aDT`�M���`ߏ_IL���B4z)�&a|�����遠oH^7n��
�Ք�O������m`���d�L���n?�F��53�A����?�שׁ�3=�᷸��V�0�L��>|�yv��7-�����,��قn">Y�b$�J�c����~�늈�U.Z�ZnO��; J��EI�Y$�dYFun�X���3�,|k�}|dA[IHI#�`��Z��HEQ|6��6O@i���,k����Dqs;;p�ს���l�'�"�s��&���4I�K=J D���v$^f���߸��8cч@�^s��E��j8��^�b%+��8�O�LBN@1?�]��b�_���ԣ���)�w5\E0����hI�4T'|�D��#�[{U,#'��b5�������l���?�� ^r�""� �AF΢�( ��n�&�u��q�kn&����t���O��`Xp$Ex�$��d����k�'�2ѭ��	Y�n��f�t3��ZI'yO�h���4�ن��>�)8MQߢr�
`�Є�q×"TE�pJcqpg]�\�#$BS�:N�x�oƷ-�� ��
�u�1�.��HC^S�o�l���\o�n�rӄ橤CMb��K�M�����tܠ3�Kl�w�X������͵�I��^a���bʘ!2{���7��|���þvn��I�W<���������G���V�gl�o]h�Vk:�����/�R$C�ݿUWKgM�%�##sh�e!ӻ�z8fK'�%wPP�h2}�w]G��0�a|�3� c��E���Rv������u���%�N�2߂��KG~��g��{+<;'RSvs� �TqՌ����M��s���?�B���@1R+��(s�N��-n���ʯ+�wD�X���Ͻ��G�����3�
�s����5'݉s����rƔ�V�h,�P3R��Q�ۻ
�~��p��Xs9��J�x]G��CxDƚ�fX��cE�����/'���}�u�W��������l��5��,fz��;����q�qvU�L\�;��:i�F�Ђ�iY�#:
w��������@��Gb��-�2��3�]�_���i�T�(yuQD=�+,j���-(С��^����񀫩pI�� t�9k���b�c#lu�	ƌ���7�p��P\\�秔iM=\�0�v��O�ԇ�"��/�2�3��
��Jy�O��dP�9�����a~ >c{�n�q�3�����3�P{|7o���ƚE�u�n��9o�	L �]�m1�-� ZN�.��{��=�M���!�g��KB��\�:�P�deZ���["�/(���1�N�"c��"t!]���l8$��>�����/_B���o�?j��]i���3�};�RT.�@��!A:�0�V<S��T&P�a<����`X�&|/{�8S��{��G��a�B��������;t�CB�y��-Kov����ʃS|��� ,)`4�Xp��w�|~<�5n�Z}�y�+�0��͔��x;�{=���t����1aY���,�'g4)�\��k�%<���& F��l���Ζ[j�a�F=��D����w�/�I?����B�G����R֨}%K!/lBm��$V�1�㞐&����\��#�p���OJ�oU���"�
R/p ������ݱʞ���$ {E$��B�w�n@7�3��cnER}&���OQ���x��ر������19C����afHq(?)��)$�~^]�`w�\�#OK=�0�S5Id纳��k���o��]#E��Z���7������[	�N��(%cY!..RH����@��Dk�I׻�m��Yπ��� �yvj�����N%TG��m�4x�1�}�	�3�.�f���JfT�,���H������,äW��S�`Vo��uo/rT
�T�ܽk���v0���d�`�Y�FJ��6��to�ƞ+i[=!�o@wP����&T�����G�s����`��W��@VĎ�U��]�K��%�X)�B˭�Qj���ZyIi:Į����1�S� ,��G������H�#�`i����6�Iܲ<^6 D�l�W�<3(f���
�'� $��6�Z�cW!2������Ox�� ��\�P�lG��<���H
��/�����К��w�ã��K�$=nR�Bx)�Ѳ�ˈk��)|�T:��A�x������j����P%�?�O�:�VN�'�9)KR�jL��Q�]G`\����8��La~&�&�L!��A�u��VFK ~���>��/<�d�m.�s���P�.Kh�(Xd��`�1�kϜ��ɥ��򅕞,M�@rA2� `��^*�	J���g�	�(�u�gj_�ǒn-�O��'���>���n��)�1j����S�������0xd�8x��e��ae�$�^l��V�5�m�\[oߝ�Rǻį���=�ҁ8��NG9P�U�b{	��$�W�����b���V�l]�Gj�a�E��[b�fI�s7.]�	��-���T�z��q�J!9j�ϔ��l�]k5q���  �E�}�&t����ԿS��*<���*��w"7���Z�{K6�F�4�u}\��@����s(`�\�:~IW)pN`k��Z���I6Ko�o�A2�y�^-��L&Qĭ�E{H�'��������
c�7`���?A�ZF���Сe����=�/�j��
dyPg�E�H���a�Aa�Ya�Y�$>Pq�,�_�(4(ܟ�57�'RRQ7�֢�}9D�o�L&�{�|��[�V�1��ɋ��=�B�y��i猶%~�4�I��͔7���Br��֏���R�4��P��I���4�{�����X���TV�q�P[��%<��hf���,ЊT|VNF����uc����11Ǉ�����]�M߭s�r��^��D�9s�-�f�Q��s���:E�.&��|+k��~��� B�".A3�����N��u���"���&��ڼ�fc��t�Rw  �HEx�$�:Ȋ�pZN_��I��7���dh���7���I�}?��(�_vǩ=-�D6��JS%�.��b�Xd��2p��Q��1<�(�������e/�-O�!��쁸���\dp����pVM'l��{Ɵ&�5���E5�&=D�g�������=S���;�U����GP���B1Ï��O9���6ԅ�@o��ۏrX�ؿY�P.�=�� ��qTXk�n�� ���r�!�M��D>rL|��]?N��l�ϳ7D����skTo�@�#�7��E�C b+v���Th�r��z)��C�ye7���-�D��#n�]����F�U4���3Zt:1��{��-��C����<����1��U4��ݑ��^<�W����i��V*uc=��}�4$/1��>�}�kl ��!^7�$5$A�r:�ȿ�W�.>��:yB(��;���PTA}�/ i��ҮI*����l�MS�*~�yFYx!�������e)%�9Fv["݁�C�&�Ӭ�bK�+O� �v��%������(�C�T#t�f�X9�D������R7�Q���ܚ�`��ؼ]�����;qPl�Xȋ^�f��>�@o]9_N���-����.ւMT��ｵ>�F����6v|�����~n�zQRS���8�m���&~
��_��Sn�=����+���C�y��{:+�~��D�;�כ��e� ByKu`�:� ���C6�CH�	U��c}kS�p���}�qBeB�]��R��ϢY�{��3n����9q�3,S��B6MTͱ(����؎-Uӣ*!N5,���lLFK��mx*|3�� �r4�����Wx2�.�~�{$#S�ԩ�6u)��}\�C��atP�p���o�&�R������	�0MLuM=��Fwfw(�5���+M4Ϥ��e����͢	�vl����&�y0�R/Ӂ:��EO|nbmC��#Sm�S?:��փ�fHKLr�b4�ꊛ;:X��]������*i<AxWr�N�(D_1���P�e���ʗa���-��1R/X��ѩ�=��ǚ9d�{{��@�T�/[�y�$E�������,��z5&ZC�12]�u�*��^=C*j~z�I_~JR��f6#*m&t��w�Y5�hO�c�b��ЏY\4DZ)���X��آ!"n���b��Ǆ�R�e'jB<D���WfԘ����3,o#�ω	䦤i���F߮�l5����M0��l���N'�.����,����k�r���	T��2q�u������'�R�Yٿ%�T��_��)�� �n�k:��-�:0ÇG��T��JG%+1I$%�sͲ���l�.�Dˢ�`��U��K�`3��p%�0j�_uT�v��&���w�q�LF��>f���a��m�=��bQ�=�GT�1�8��.-(�e�%�XtG�b@u��4�^���1e�����e�N��C�n�v��b ����l
����9*������#��A��p<�Jo��q�#�Ϡ��C)�,�Q��pF5ܺ�X�-�9�P��Rc�����+B��#/���D�P�ak��Y��L,��a}�_n#Ku�3�K�'���*���,)�����,ELx���E�g�j!47���NŃ(Hq?SG�Ͼ0.͈1�{G�璣<�ۍca�>�.�?5��Qi��М�}/�OZ���;"�
RGݏ-�c���h��Xz5�֌�j�;g�Vf���f:�nW���
�-$Ipy�^�c��vb)���aפ���T\�T�7�9�j�[��-r��q��-����7���615E���%�ZST8D�^TX��h��a�3��_L'� L-�q�0�� ��\���g��!U�y,�,~w�2�(]8W��;�@�~�I��lz����I�[�x5�:uW�Zl�X|U����c�ܥL��b*�P=*�DDp���ֳ�Q����>������ C}:��Z�`��bMX����zެ%�j8퐾��"���gyfl�9�'J�ꖙ���}���*� 8�]&:Nk����4#���K��1>��S>�����lf)ь܄t��mr˟?VS
�)�kWJ�K�
k���s�:�nm�z)sIw��6�s���oo�$����nɀ��4PqR��K��2��ӞJ]%^�p� �~�_�/�u�"X h�@Aؾ��bl�t��w�1��%�S�U:/�=Ic��)���Pz���y��C�"8a?<w_��C�@�2�g���b���� p�*��L�*9�as؟�\�7�������J,�˹���^�?P��n��_�����޸���gI�*��~
���9��������u�ٜ�)��Q��vh�W�4���>M<�۾C�⮢���#��KgM� <kU}B��A��x�>>�@����NV��eY'�)��$h���a�q�1(&+E��������NCV��z�qӧǩ�~]����sl��1����_}���J�W3�3��>)l��f�QG
'k�{����+�=��}�FQ����Ⱥ�Tw��vMF��͞>�%V��e��V:,�쏐;!#�W�,�:�c����keK�ybv��aR��T!����uB�,�a3?{X�8U�~�(�ƒ��3Oy����4e�a��S�bHؐw��y��FR��ˍԲP�/�e�)6s_�����;�U$f�J��RO�|a�0@�;�����I�P�1����u�,�nX��_�N�0�& d�c�w�d�i��_ Jr�3��&�	�>�'�=���֭qVF���6�`±��=:q��@���7X2���Gŉ�]>ĳUZ�<�=� N�� ��bH����rȒ��D��l��"@N�kf���Bb4(�	o�i;X=���f���z�]�Ӎ�H1�}©R�
�����H'�7��'	܁��j�����Tf\Op5��t܃�N�a3��Nu�-iB���E��
�!Wo�^&��1<���������3�(�չ'�B3n�K�A���a��E� �����q��W=v��_�'����]0�cP���m�H�؃dC����\��b������zv�g}L3f�F�f�������7���=������8eXiP�s��[�HL=����>DoYB��}(K�ـ�UUkVs�,y͇�^lR=*
:��mX>t$�WM��et{6����|��n��a���a)�5)���(8�~!2T��=E�) i��^&[��W4;WT7�t7#:"}�eK%60e�:�-����M�+�/�h��ʚ�r7+ׄ�k����z�;6��p`#�ڣ����m2�,x|��L���\ml96~�x-�h�&
���_M�� �mA���`���2[M����rdR�z�r1w�w/fT��.\5�Oc�^�.bfIR�y6w0wXQ���MNꩼ���weY�E�,�jq,%�f6�ΚǇ�v$R�h������q��H]�c�Hb2x�/���G$iE�߲M5o��8ɋ��Z.��`A����S1v����W_!��ȼW;�>��e���)�|�B}���
H�%���r!�� �W%�h���x)U����TV��`U��4$�<Ί���+	�
��J�`��M�r�*��]�H�0L�V�N!>�J]2C�od;��㤇`p��l�y�>��=U�]��BZ���, ��n���R��(� (�p!cb.�#�?�y	��Zr����?���z:D��ǃ��Z�2��o����1��i΄α���9��v~U��2�ݟRpw�E�M<L�����z:WTgh�Z�Pl\��ÂE;gs�F�um�m��!h?^����uճ�1�
��`d;��VC���0y�Bbt�!� ��;W,p�˗� �6��%#W��!�j�	��3����茸���^1U�bS���귈|�j��������G��u ^Y�G-�8��x].Xj��	��M�N۳�޻��׍�q��&���IFD~��	�o�3.�������ί[K���V��*uf�'瀄��r1�TF%��{m��9�لF�-�m��5c�9���T��d?��J-�3���AMLu^�7�9h�znqG���u�P����C���ha8;x��f5�m�u��L�/��EDK�d�Nr?���m ?�ifJ�mHC��>�;H��JH��°1����Ƹ�.`'����C��Q�S1����޼B�wm��@�&���w����ňRtRI�R@TR�2(�d���Ō~w��Rt�,�
��¡<A�M�{���Q�q��S�c��n���.�N���]+�to�I�E�R�JS]�=�d*��Q����;L����~@�9#Qv[^��|��!Iu�v�;f�з�q~�q]-����R�w�{�1�L���ϱW�] 4���UɚH/x�e�n����R�
�G�3������?���W�6B�{~g�����E�7]�5�l[p}��k�%�&uX��
�AX&&1�Pb_ʢ&�w{I#��I�A��ޕz&q�b�����M�!4G�~9�p�X�@�F�A�DbS쌔�w��&��\�$d���|JͷI��ۀQ Zcjq[F'�g@�"�:n���=���7t�mz��J�W��	�� ��mC|X�n"�ꈃ��G��Hz���VR�iڀ>z@�^�/Cd���
[��t0�N1�S�^Ӈ��Y�K�,���_w�0�����;�N$�����\Y�Q�E�������@���e���h���7�onؼ�!S��K��Z{}�_�`9p�I�7�ZY��ɠ�e2.3:\� +﬌��)<'��)H��L'��[�T��Z�)/���˷*���C��V�QU-�J���^9G[@��*�E6�C������q1�BK˭
|��}�mL�Lzc�0I\�,�y�lGm���\u�1 ���V���>X#�r��ۡ?�xI�0���*�/<|F���8�+�&�28-�!��}x�ɧ�0�9"T�d^N��F]����x�tW�u��*{��� ��	�$��4SBpAw����D&����	�ĥ����rE�����B�%���������K\tNclKPB�e�:��վ�2/*��w����޸F
�P9
D�Ć
�@�tM`���ʌpZϰ��s�y�u<�,�X�"��.�U&t�ա%�:�d��)�k� cQ�9�Q���$�5?�h��^\R #ʞ	%���n�⯍^Y��Ta��)�Bۿod���� ��۟�ܬǵ�P��_ɧ�(o��^�=�q`��iEuF}��͡��"G�eP��w�����VrN�X�ۜ���')��܊��?V\�����j8w��k}	�1Y9�׹f���r��7ճ�gը׉��`��?���ǳ��)���h'<^1h�pM��}�U�a}�I��6�!�HC!=��+�:e@������!9��:����^�A˕��Z&2����,N�tV�[Oͳ��Hp,�fh�dK7�O�f�7@�Ciҿ���O��͌��d~���:}��@��ן6�3��ӽ�V�c%�H�C;OV���-�T`$��J�����aul�M+��c�OP[��*��H�AiO�	�K4�߉�fT����i��&��M�7ؘˬ�Bd��H�$�a*�&/��t��tw��D�ˮ,	�Hq�R#Å`iu��AK�g�/51%���.3ïB�<�#_�t�4Xlع� (*��GkfM�����	�lCX��t�4�����(B��^ڛ��T<V�q
��;<Yj(뽘���
�#�д�|�Frw���xlȺe�p���'���hf�$7�����>�:�u�U�wP1���ؕ'��!G�	��R�k����������tV�8�4�{:�*S��"N܈t�굦'o���,/�՚T]���ᭋA�:Y��2��_\1o��0����~��;
\��oVH��pN�vܓg#��s�6�L�S��2|�Hh�m��d��KHc��~g�r֊���`|ߴ��A�Z�p�B��٠��]l����RN7n-q��U��T�;��"d�/�t��� ��?��U�>��3&�;�8���eh�̌�m�F ����2noD۳�Ho1\ 䌝=|�kN�w0��'�B>x��S�[�&���g^ �������Wf�T������b(��"ʥ�
8Y��]a�t�����AU�2�r%֤�Z���k������k�L���G��v�,�:��Ԇ|�T��Í7����7@}9����)m��cԩ����⎑������V�~�~w.k^f6G����y�������Lq������=\q��T�N�G���݈�9��A�?$Y�uX!֑y�P�'�R��#IS�\��/�!3�h��2��7Фd+�aw��[��=V��9 g�oQ���5�_�Ul���5��ɬ�{���I�n8��6�Y���]��f��^������r�_O�=�d�)G�����h Q[��+T�b��V$�.j��)&tg�e�]	�F��1gX��7yi�^��W�^s�߆!y�\����	ŝ�Vu�
�\U����}����rØz)�×J���'A����ps�)� #g!aݒH�;����Q�&u��\
�^#�;�^�g�'q�RA�gU�F�K����:� !,۽�L�yeZs�������h]�8s��J�N�zN�$f�k?ZW5����JwC�i(����K!����h�ҮU�5���f�}	�23
/���zJz�]͝+"��X��D�S�[��W���[�Yr�v�H��+��Ȝת̭�f�����}b�5��>b�33�|_r�h�2U�L����P6���]p�D/��P�r�=.x�#����m�׎h��]! (��;�į[eF��.�1�Vs]C%�X��=V�/{�L��Q�Ƨ��ݡ��CG�i�.7�]����'���ZT�TOJ3r�RxwZl�c]C�Dn؆ �#l1��_[�m�{�5$��N��W�B-E�g��Zѐ�E~A�.6��џ���2��� 8N#��C�� 
���WAVb�)4D���x��q��1F��*-�!h���=�>\C�]�qa1;���x��@ޏ@f�*��Y��L��=��,�4FޛUԏ~#��iv�q� 6z���1�+���x��(M��z���r�4�8R����@T�� 0��1�|����bS%�N1�˅D��.����;5V�)��@d>��;>�g���a�ʘ�!(���d���R���pV����	1����v��dN�bj��)[��?�1}����L��bL4gꌮ�L~e�r���:(h�{Y�����u�
*��
��#�!:`?�7��T֫���4Y&y�f��9t�ef)à��,��\�|s�~Y�~�����1{�V���[�!�tC ��U}v��WL�3u:d�W�3U�9$��)?9/�(L��ɫz������q{�3��GvƂ���j#�!�A���Q�B��QScp1u�1߯=�B���?Mf[�#�d`�#g��(|TB0S7Ӧ!6s쑑���� :@i���l5�C��m��\	8���U� �J���E�c���/���nu����<��l�H�*�����J�Lg����$;���P��e9�Ȕ�*�w #��l�����Rj������a�p�u��ڍ��G���u�6��B}�ҜЬsq����+���A�}����8�j�t֌Uǁߘ�&�Kq�>]�J)�TƋ���"��ˉ�H����n^�sՉ��̷�t�����W
��>��i���%"�q�v1�|�
W&��~ޮn_��Q+6]�1��'Tc�*�@[B6��`/��vI*�.��C���vu�e!����	�8�FMyr�-�3�(SbRM#t�"D7'M��6%y!��%#�$v�� C[��iV)Ǫ�8�X�o����<����w[?CBq� ��a�˾�����RF/���R����ha%�4&��r�z|����0�I��z^��'"��pޫ��1�qc��o2]�����W�+��!+F��P\`�l����Y���H�����_9��}p��`_���+ݏQt3ɵ���hsd���:u�)G�6��p�dD�׬쭱�����W�(��� b`��_��L1/r2�O��z��r	e�PZs�#Of��z4��B�5`S��ʏ��YO�av��ǂVn���uu���h��z�4:��3�gpjO�^�0��RK74ԑmD(� �KU���]�d���S`]'.����ڸ���z�$��J#�xyI���|���(���8YEP0�Rd�7*ޣ�h�~�<�dC.��.��btje�}�[�|of��ʹ��P�-���������
�h�n����t�<%~�����<�V>v�6��o~Ųw�.r;����eދ��~��1AT�5�UwF�hi�Ӊ\�������q���>-u�'|#+�j�ז�u���|;�	�Q)>s���PbNH=<�w
 ��8 �=����N����w��l�}����x�(�/�rr����B���.���#����+.)P��R�Ι��GM�R>��^�ʫ#�����C����Tz��l#+�s,d5U����D�y�tۋ��W�Em��&�7��4r�/T7|���R�-��_�P��i��4f��)�4A̟B6�#��:�
8�d�F�����,�6���Z-��Q3��@���W�L]��J�i
�qY�JS�Q��a���l���pj�(��0�r7�5\�#���� �O�{��!vgu,f7�}>E�zPU�ݗ�ӵ[��t�j�6k�N��0}l�;M���6%Kڊ݋��-�s��G��s�%-6��e�w�ҧQ q�����	hp���`�Y�<s�p�[�D���K+v��D��4���x�R�ʱ�>_^|���m0���@a���x��W?�͋���Y��*��8
f�q�4����F�����"�d���Tr��o��m:��r��r�g�s��n�����>\���y~n�~�ȈXT�W^H�C;E�^�uy�|~�K]���6ؔ��a��'�:N���w�U�Ҝ�*�.��<BGt�wiчIS�FM[�Ҕ=2��7�+\�E��*�CD\%�6�`��P�`bHv����@����ͭ7��B�`�>s�^��4Gm�I��ͺo*̾͂m�*�r-Ţ�G)7�T�����CQ�'�J?ZFa�\��Q8Cx.P)VC	I�w�г:�Hx�{
�{=��T�ˎV�X���'�F��A� �}݁��%�J��U&m�B9r�&�wگ��
{7��Z�)z�~�qq�I%��)�[|+�+:zk4m�e\��`������� �Ram�¨�������@�h"[��bM ~�TG�8I?z��Y����/�UI;�nӠPB�S��+z�qT��tԢ"�"����;��@D�vQW�����)���p�Uj�ͳ����^f���:��>�?~�i�n�K�\%�����N����;4� �`$/�,;�nh��"����Z��s�v0z���u���������)�N�:@�n�օ��Pkq��_��g�7�Ì7��k݇&7W��k_xmv4����<�orx�UZ��w��w�r+�ԇ&����m��c�L��AA�.��9�����i:�J�u�q���ټp$��+딞������by����Rl�Q-���H�f�슐����K����t蒰7��^^�?��׫5\����EX � ��h5ď,��?&G]�w����^կ<v� ���3/�j���lQ`wvZ}�>��ubL�}���/	�e^WiAdko��A���v�K_lW��ʊZ�MxZ6q�7���>o��U:(�7G#�H�6��aN�H��l��۟Kuws��:�#+���-��J3.���v-	���PBQ��Y�y��=ң>���i���F��_#x�ea�g�A߂k���r�.�������˫�@#�tZ��7����Ϲ�^�Cs���G��g��+��ȝ�*G�*n8���S��4o���/1�5ƕ�+�H��$�@���|#�,�gTv�W�)��(aq��햓��yvn���%
��
�� 'Ϧ�%e�@�����}TP���}�Xt�)��C<-���po�>��9��)lT� ���4���!�E7����-m|���Daĉ�sܸ����3]*���XG�o8��� �x�1k����X���91��m���9��(�kUYӈB��"wxL��Z�w�@Y�;��m�UnS�R���Jg������K\��\�;Du���aN49M|���%�vhr�_5�E\G��-1�o��$vUMS'���`6G�F8�--��]��1[���{[*����mN�?���cZ�YB���,�����x��5m�ZH�'O(R@�wN/�QU�,�&�%��3*������"�<n+�f�h9��B�)%�4�R%�y�V+�3�>�=J���?>�ʚ����*?ǁ�o,�:$z�e	����'�/����M�	�P9�겏�� ��e����pʅ�@'M־�mc����������w$��*��q�7G�^3�m`1^#ݕ�*�k�j^�@�H[Q |��"��L{1�yDᰗ��<�F�0�@`8��Ƴ�	J�8��ZZڍy�1��������#�{�C�9c��ra��\�R	�=h]fX��+�����̅�+MA�?D��v�E����@Fn���n��C�c�(�$;��&nL+�Ψ�}a��O��<]�u:4QY#aQ=8�Ft	q�4������ґJ�M�_���B	f���2�Xu��u�JH�R�?*8Z�T��S(8�bZbxG?���uv�F�r���ؒ�x��s�
�����=���.�G�7�Ī�]�?�8�]�@��a��خ��GN߲y�['�|��B���vs[�y�̮���e;X���Ik�.�__&��BV����xk�h��Tkf���F�ζ��^j�ghʡ����,8�8�/ �Yv^v'��]x$6�d�j)�<]i|:��U��9�e�<�a��V�B��� �m���2��(��79��Y����?�?}���G�um���gO ��,�,]䄋���R�U���:�j-SJ�Z��/�KT;dXPƏx���b��@�F#t�%�?��z���r<4F��>5LIEQ�U���í<tmlԏ8��K��j�)�6���h,����A#��e�� U��g�Q���.�ix��or
��N�0�4e�A�����%���)\3!H�P[+C3	3����1$���,�����U(�ў�p�����H��HC�<��}�-�=POZ-߄��au�����k;Zx�ر�mu1V$��O�~�h�;h��&99�%�%-�ʁ������Q�=�������x�Ԃ��.Z֥�GV�@���\�d.�GOm� ����_�����BU3�0��P�	z$N����zc|"G6�oҬ���q��_�L�6a�7���!MsO����Pf$y c�j>�ݡF�V��9��jɰ X$�8��?g&�f���\E�٦+.�lt�ʠ��6Ήi�u
����ՋDIf���a�Z֋ �t�v` &Eȸ��a���Dҽ=(�_������m>����<��m����+LIƒ�	�\���2�rp���-K�d(ݤ���gږ�� O����_wnY�}���� �]���wM�u-"����n����Zx,��x��Ӹ�bl�J��Ip�~��I�W��{}�pO˥`�]�vݽ{����&D��ܿT �)
��ʇp�X./4�M���Z�g2��5F�?�A�>.��]�������^��*��['y����p ��Nu�u�a5Mݴm��T�*o���:R�r~#4}� 5sf~��]�o�ai�/�Dq�| *��M���Dy�k�:�I���`��M��b� r��Y������<���?|�VĂ�y6�e�j�l_b8p�$#�g����4�Rw�Q��Um�K�\�m����x���a:Dլ�cXFf��p�,)D�4��ӋJ��K�;��"��Ru���:R��w�߅Ql�'�h�;��趜�i �] o1\4�aY�u-{&�mլ�X!Q#~���lko��@��p3vߘ�8����AĵC�Qřu�Gvao�%5�=�@�9��J=�9�-�������!f�
S���@���P�$�m����ٟ��l�cAs�O0��V,k��9k�U��;�"� ד6�I�X�j��l'n�>��	�7�rQ�����g��XU�Oۘ!�P�of8�|=%d���X�m�u�V��Ŭ͋*�ec:�3ڠdW��,6r�X��K68�%��t�c7�R���e��V��+Cm_�v8����P�G��+׶s��;���J)���ڑ�V���"4L$�Y�/����%i )�������%V�����Km����ST��=�G�
��ܕB����������X��� ����@>�f����-�=A�Q�<����Ղ&��/���p	զj��QPsϹŀ���S�{�-r�.
9���U��?ؿ:�-����Z�3o��<S+n\^���x.���{�ể��uC�<��aTx�.�\
�zI�\O<�"K�T�\��W�$���0,�yZ�%3�����|��w��H\P��O��_���^���+�	#��0Y�f�=�&�aL���G�.GZ$�|#�c(�/<��$B\���s�@(O(C��c�͊��&�J_����L�Ƽ^<�bD�6p�������
����@a�+�89��*]�ߊ��RZ�ӺS���B��:���X��,ՂR�����#�ޑ��^yu�N�#q�\z����`gN����G��&^(8�������]��[2�)bY��M{�}g�'��s��+��:n�:Q~��@
#��Kģ�95L��*���ѵmΩʇ��$k�b�կ����v�q�>�WÉF�B��T?h�m5?�>F4)(Ͼ&��x5�ptcʖK-�p<��`uf����P1�Ee�����M�J��[J����dki�llQQ��C0�BO��{p��X�nЊҔ�2��L�Rr�B(���6��I�n5�� j��Зz��������G��(X�{E�]=s����5*�#馶�����t�Z}n�)^0��P0J_0�p��eY�8�E��ʩnL���bޖ����jH�E�i��I��[XN1c;zWf��w3��k%�=;�6�k4���gҞ��=?��N��F2�ۿOn'z�nE��d�w
�,uS Z�qhMF�~�Q�g�	q�X�S/���� ���ZYd�@H"7c馝�g�p~��xB�|�6����V��t�$��~��xcZb������$��[ǯHH���mսA��fΑ���^7���i���F߆r0)�?3�Oϋ��Ѫ�>uͦ�{O�!�sx�G*�� ��ֺZ�������692^Ԙ��;�80Ϲ�Z�H��!�
���ܵ*`a�5�D)�[.�iEsN/t���J;�6W+��Y�T�?ݔz��b�]�X�I�D3ȵSa���b��h@�!�y�q��f/�Ĕ.%u-H�Z��*�@UqAb:E���Z�`�� 'U���#G�&��=_���k2��E�N��l�"J��
 t��T�`��Vy��YYd᎗�X B��'� Y��Vr�'�g��Z�k��8��U���Re��h^��x�T�"Q�}�x��+IA{�MX�trj��]�%������:u$��|��[}��O)_�'�q��i��z�@�X���U#�Y9��/^���T�V�6�;=zل) �[l�3\��Y����C��'��)/S]Y.m�fN=�2ă3`K� �^� �����L?�b>��r� ���H����ܸ��؉��wb�o9�� �^g����3na����ZL��:b'M-׵�`����1�����{��4/�?#�V�4OZ8��4z%�A�V��I��F��-��'����H�gK���v�`��{�6	�V�a�m�\�Q����)Djq��e�Sr�g�7�ҍ����jk��R�؛S�1|�9 "s��
���h�!c�q��xԵ�h���K\����#O���R��`�*���%n�k3j"K��>����
�+,���ʿ"��I�����>��x$2M��{�6��:��=%爽��۔"��iw�$ϙ��~��ģ'{ea=�*��Yկ|�<sy��6x�1b����4]+u��C���:-ޭ�uc�؂��	�=�.� )&��d8��T�4����z��еΘl�[\�u���f�L0Q������9�u��=�ҡ���4�V7���K�����[sr��.M�g�qzW��3�8lL���~E"�R.���ՉI�-���N�#�� �I�N�� �	�����\Irrd�ɶWk�gWƝ,Ze�Ź���5=�q�1�zf$�/��v��v5S= ���q r�j�E��bQ���*i|�!�s	�x�U�'��)�9(����@!�h���С����B�t̞<��1,_����;ѧ��j�"\~Q��HܬW5G��>s1c[�bo0Ң���:��w�o��pʿ�I�^� ���`��u�D���Ƙ�o����,.���AN�F���P��JvLX�i�ϡ�_��JYyas"�օ��b�n�P�R��r���ie9js��dIOf�e���&X��%�ٖ��o-%�#do�N5��o��'N�4ό�	E*�q�v��"�@�ta�(B����IN�9i($�şF�yܖ'H�/��������z�4�.��\@�����g��7Ѕ�k1p�=�Ա��N�q� Du]�jw�a�N�:?Δ������[�`��%l9L�I�8x��V�x�r�P�:@���Ls�6&��\9���ʞ�Po/l��j��T��;��[���u�D�wO�i�Kӷшk���AR)Ԇwo��~x��B	�iʦ	�3����<�;�����bub����u�̇�5��ק�
%>1.>�CO�O	�/�Ո����S:��RJ(��'J
Vw/#�~��݈�cRt�9^a�o��4�Rv1cd4�#o��|��(�<[@!�yڛF;	�=KIsa!+(e7�����Jr���(~�,l�\�<:d�5I��h��XT*��1����'����s�w����W
ڑ�p:��f?ܾ�KKC�D�^2;�ѫ�v5��m�Q��:(}J<�f�[>Pw���Eo�xx�S�=�]��p�i��5��?�Ɋp�d&ϺWe���+�<��Q�N�cMY�� �[��;��r�@G�/��6]?�G@B%S����@+��`��|�I�d3�<�jDHc�!o��z�Zt��i];�r���P�=��N����]W|�. �(�9ʌ�]��M�_3��͜SiPFM���]�0�VL�hfc�o@������y%ւ�^P�c���@P��]���[�S����^TLՙy�����nA>���I����&)�C���H!f$WH������8��Q��a�@�0+L�#��Ԓu�o0,Á�T����#G����Y�a����I��BA�jܥ��\s �K����� ��6"y�����4�E����t���W���+p�1�J�&���Y����F��T��.cj�����g��8�]���"!�ja�{%= ��0[�ɥIc��Y9�2'��ML�w^&�Z�[�F,��}+�tS�
�ĕ8v��j�a�dD�A��2�|`�2]�v"R���a��p�f�Moŏ[pY1�� �-�$	���1�3�zq��xJ?��`�hށ�9�ՠpo�@sv�Tӎ�1���R`ܧ���i��'��YF���&5=<z�����P�5�y��L�Fo����r�����廳�M���Y�z���"�
,I�΁㊛w�����(0La(\�$F�{�3ִX�h'X4gd�z�I�[؜�([a���1벇W��7)F�E���[���4\�m��tY46����D�էlm�^<g��Z��i�`���񺦓������&�TR��Jp���5J��|;��E\�%, ��x�|D�mD��f�*{�L���Cd	o��;�u��3r'���E�p�'ZV��A�m�s
[�<�p�E�3��m7�gw�s݀l������E�`Ի~�7����~2��{5��i@*�ׄB,/N�3_6�Gh��2�O�=|V���PygEk$�������nP�����������`�oA]=p����vf*U��Ovmv3�z�6sM��4����F���N�l����sc�41���Z�m`Y|�H\����[�c/�M�	sq�`C��ZDW�����'���>ʺS<X��)��^¶��p�xyRӞ!�j�����~x��>EC�{ѝ��	Al���l�b�@R�̓Շ2[*��*lđIH.ëѡ�A;]@��;� ިx�F��E�*{k�0��KTx���f#�3��3�K�� 3�e��A8'�~���O2���[/,�c�z�}K���)����!�9�Y��Mrp� �!l�$������]N�}��m����
�A�cATƕ��U�(����.�vJ+LФ���0��Pр��VDDh1� ��́����f���Z!�҂�qeW�[=)�uT��V��]��Un���D�s��6$��qx���U���Q�KiB Y�W���S�Wcߕ�@ӱͱ'l�h������O�P��MX��z\����V�`  ��$��[�������~౪Y^{W����݂��zՕ/^0��
0�"5��@��G���T�
bH�;������� �j�n�J=�@E����a�N�����+�J�� >�ͩ>O�i4`� rw�E�5*��#a{�]v�"�����+��l
���kM��Eف�|�;��PưS�~�T��\��"���0w�ɗl�c,�}4�TvH�%�n�{4Q��8��o��M���&�d4"�q�p��I�2��6 =vk��]��lPe�`��;��V�`�+\Bʥ�o���l�&QZ(����:`�>|�oF7�zU���i*l���L$���b�2�"i
��,�H�k����9�I��K����XY&b�<���"����u(m�O�!p
�j�olIN���V���}1u*�:G,�����e<���W�^�$��^��N��
�M_7;*� ��Co_<��K�S�֎߅M���$�t�&l�7���]gw��7��T�o��s���&��P�~�@<uN�!��
ɑ����qQ
]��.��̣�>r��`W�;{�n�T['�CY�_
�=I���I	jNs��o�N1�ʏr6m�!�Ǟ^W�;����=|�j����N�JLpD��g��v���x�9x��O��S��{p!���)e>0�#�����V]Ka�PہB��S��?d�#��!\��|����I�X����%Ʀ���(}��#��{�t����
z.��G���+K��������t��̮��qY��>(�@�� G@oo�z�gz�۩�>]����~!�k'7�UI�.<��U, @���vE�`�goM�T�N���������S����qi�����˴'|��Э^t��p(^@����F��J�D��%�������(�}�{CDC������Ձ���j(l���ˋ/����";:�|JK��4����2y�/'tV��ͺݨ$́H��������o��u�46`���ޗf].��3-�(4����Α������򘋀x�T;˹� :v�KE��̼�위MS!#��#��8./g���`hGXc��"�_�k��������yq����-^�%C�Q��,4+�����&�&���-v�()gt)���"0@0>��%����z�ڵj�t�h����d��|��	�Y١a ˢ6�_f�U@/�boP����=���Ȣ�wb�G�F�<�G�c��ҬZ����w��[,Z�z z(*�MY̘�o�ٙ	�С2N>b�j�}YЧq����Iܑ���J��>Y�gLD�&F��H�K�|���ռ�QY���4�C5���\�%.OΝ�z\O��pc:J|l9�ϥ�Z��0%`<K�6�;$5�Ԋ��r0`I�>8\Ь����:*���Tb��`s@μ��
#2�./��]NH��9rLI����v�F�hb�$�f��@o��4��r7���6Q���<^�1Lт9ۏ��e�dY��8���t�`]\v�Sf��D�!V/=��;���"���[f�8�w�W�e��M즘�4*� )4����������	�L��+F��1�iRw.�̬�ر�4�*��.�zm�)��0��}����g�H��fh�
������Zh����O�k���ؙ�f�5�K�]8����-o�޷������}L2��H�#�Ӂ8������d��^��J@}T]��X����U)l"$u ��xz?�3	����ֆ&���G�7u5�?+zO%�h��t���iMz&��z!�Zt)���B<�B���|,>��pwU����&x��(3��i��"�c	��R9c0���v	!��.�JB�P���b�#�)��HC�����q�݅�Iu4��r���^�>�܅�n��.���� c��\~��Z_�`�z�u�OU��sF��� 
H>��,#z*�sЎ����,�BXπ�z$���2L��ۭP��{<�{
�-��)�J�S�N��7�)�I�O�U{�#yC��H�<��c.����)�z4��^Or��2�.z�tWFV��
�������`��SE�/!�b��wA�g�������0�w�Wn+i[��d�F�!%��XbQ��k�y}�"����N�4���)�t��H�~������<�r�ΟN�����E:���E�t���c���\���4���T�����K��Vn�ױQ�"!`�@+�А��Z�K������=�X���j&�DX��܅���m��i���MFTg�4�y�aֵ��l]�)UfXl�4_���a�ʣyY㶲1�3<��{	��D �R��SC.���u��HU5 �<� �N��1�l�Ѭ�g	��Ae���t9��B�dpk������f�޶d�`�O�BA���Q�.���'���9�j�0�uY���i��=	o�W�ː0�-���
g�p�� ��]o�ERHb���p2���I�&��]�x�����m�8w:�C�K���V�0��0�I�:NQ����b�l�u0	��Q�I�Ib
uо���g�,y�YX���]����3頻�.�ʞ=��
',����m���e'V�8NKɹ�t���)�h)W~�ʴH%���&��-tTA�njW*�|�!:�q1W}F�T�8�D��#�J	 g v;K�����z��c檠��� E���u�!!PU5������#��t�R�j��f��̈́*(�XH��[vR�&nŪ��ςx0,�=_N���@(%���Չ��z�Ʀ��<�x��z�����ȮX~�jVӈ��|�t��~����Ȃ�֞1*�_'����C��}��p)�����#��<�_��#~�%�w�t��r%�$Tm$���T�����pv����vMF݌V�0{_�>NDR���P~��G{&'_]m����ˆ),?�A�͔[H�V�fe ,*n|�"#���Iq%*�_T��Yo-f�	~dH,�PL�d�ⳡv<%%c ����o:�g!�C;��<��J�S�R�5B:�	��L��V����F�E�]�k�׋�n��9LAu�ꤙ�Xlm�
Qץ"���0����\�W},�G����@��0Q"��h>9�C,��eDM��,������Ì����ՙ�ϣj�����N�
��O��w3�Q{ԧ&��0u�0���!&<��0�4�ѹp7q�ol0B�$����ۘ%\47ؼ�r*Kx��x�1J���6<���-y3u�����ӵ��P�^otZ+��
?	^�f�y�rz�F׵���+~E�$Z}���̳�-,�TO���Y�R�V��r���N��ҍ�9Cx��ttv�@��S�dC�R+�։������m��޸�J67S���GX��＾�W�fr�US�N��3��-bA�gP]�X�P>���y���~�l��̰�����:R�����AppE�ɚ8��OpB�P`�=��W�*����i�cߠ4�Ғ��kI����pqŗ'�*GvPp!"O��/!9� �'�7��n��JI���aS֮��pBn����Ɓӗ-������},kc2�y9�F������'������I��n��ƾj���.�$����A��S�Kyj��J+s�xFyaQ�-Ya�4��	�йY��e��` �(�ڗ�,�r9�4otܧ�<:��@ָ�:��ݜ���Q\���r9�Q7=�v��ζ=��o�����l!�gy�!�CY�Q|�V�z��v�],�@�Hx��{g�8&*�K�g�"�п;��`����}�������$�@�ΐ���F�ƴRH���E���+��w��f�E�"kj�_�n4%4��`�Ls�u6E��K;�ˌx I��X�`�g�k[-�22�Z���q���Wg���
�8z���,g>�*00ɘ� Q�9��U��ޑ�x����U7�
��K2Է9���SP��t�(��	�#X��<�9}(��P�V�I
���h�<�˞[�����oH�9�s�M�vݛ�X�G�7dwa�;VT�PW������C4V�!�Lbs"�����P��}������]�(��H�hÌX���_'��l��;��=+w��'���l&5�4۠'����7~ذ���g�ȇ0�����s�F^4��M�������Z� �o���Wc%2�6f�zO�f��w� ���bW| �ϡ��>R|���ٹ�J�'~�_���	Ϯi����%P:��a5�Ќݏ=W�=S'iYd���F����	aӊ��b�b{��7Ⱥ:(
C����u{�
ݵ��C���h]^Jc����� �IC��|7�ަ����{�����^ǟ�Y�#�g|�{=/��,F��}��m<$�O�j�9�e!�9�u���o���stl�Ԝ]�Ftp��L\��6���w���!��8C~��`A~�����h��c���Y>����v,��8�پ�r��EsN��P�bm���:��5�a��=YD��a�i<�F���$�Ҽ��p�t�b��E����xϚ=o�0��d��c���4F���*� @��y>���V2�4�Z��7��C�Z�%[�P��Ee�U{u����0}&bq���ѭ��ZM����\wy�_ Ny�q����փ��F%X:9(��б�#֭}�=�������ц�{��Έ���;�Ӎ�D�'��#j?�(����9a)�LS��8��-M&�lrmkP��)|(a���\���7��du�'^CmԞô�0f
/�w��"��Ѱ�C��j�͏4G����ʥĮ�+u��De�)-�%���W ��G���`ecAә�v���$�?�i^e.���}7�/fI��P�M�r�|�IT�$v�5�4|5�|����4�Ӆ*� ����.�"R+Oi*�:��j#&E�o��s��_�J����t��W�C= )b�m"Y렔�[봧4�O����s�ay���D�$�#�[v��p�z��5��o���QR�w�`j��\r��u���OD�o~�ow;;��h���U(�K�~4�^`PHG��Z���Э�镣2��I�x��l�l\�|3mU5ڶi�0�h�CË�"mS���*w*yHVC�` �~#k�X;hy�x@��V���2��&Yok�}�5^�ƿ��e9{j�������BJ5��d�}7�wkk�~�j���?_S�Uuڰ?��@�CWT�0���F�v��F����7sm�S͞Ƿ4 �2�֊�i�(�VW�b�����;Wyv2�hּED��n��Sf)0}�@�*9 �x����5{%�����n��/;v&:Yps�Ā�(6,��\bB��3(�)_<��A���G-��_�y�&vn6���U%��x{	'gK�;��a�\�F�}��dY-����.���	L�<� 6uj�Y�O���6~�'ߤE�uD���b��[��Y�xà�`��0�����lkh���;��w \��.`���G��j�>-L�ݡ����&�ew 5I��-3S�� ��o搞�<��B5%�b퇷�'[7�l���v��m�|g0/*����5}؏'h?=����b"w�e�+jt�2,�u���J3ү=��F��on|�)<+��9t����O��qP��}�ڟ��ܐL�Sr[J�@ޏ���s=����V��ٛE��P`�J��=Oeԋ��a8��c����Z`C��Ia�E��׫>u|w�6���6V`����塥e��b�	!��86��Y`��J����/�wT\Z���3~m��х
��5~ż����nA���p�{�o�͚�l��!���٠c�r�.���f���	%Qb�q�oY.�H��-{�+v�Y���A/)��� �e1Mj�E�M��'������r���3�����l��1��\�-zQ�j��Ϥ�n����Q��R��������Q>!uC���#���y����¤��qz����˓��-��9.�J������r��9�~�P�^<r���)0��U����"����L�@��p��9���~��Q5f�w�����_h���F���	k���H=��I:��`ݰ�	����k��5�%N0gy��l��lB�������)U��
~a2�?jWp�?79	]PWbᕡrV���.
һ!��
��R�3<,�:nO4]�r(17Զ&4gc+q9z; h������3g�����p	//�~aٸ������|�h�����-�&n��oa��	�*,V6�@t��U3����	��}:d	`�U��N[������Y�@��M:V�#ҟ��o{OrɮG6���P��ygՅ #U���%��d��R&x��y��W&�qt8d������0�j�]�et�42����X��D����`^�����k�����,���db���_uI+�-��csT�P����'8d!�qv6���?.��C�!ϋ�v��H<��:XbT��.��~��0+����i���߇��e2-].�6W)_;vSh�$6jZ��m�>�&+#�N��	��y�+w����9���=c:�ߌ��>!��'9zUv��4�L���%f��te<��h3�W�k[� �w{�I���}V-�Rultw]�J6��%E�����w
k�m>U��C3�%3��ጘI�������B�1;������4�՘C|�i��g71K0�	<]�3����������фd�M�*��IX�^����td��%�O|�o��2Ih滊h)(f���͑\u�Q�(�9�G�!aH�|��Is4������ښ�����rt�s
�u���K&�5'd e�/.�-x���g �����o����+�CIU�e��pX=^��1���+A%	H��~��ȫ6m2�Q��xp�����S�������9�L��-"�G�С��p��$�����	(�)E�p�#B��[�����y4�:>�K(�P(��k���]sY��sc8�ɽU�<�ܰ!�7�O�j���9^��C�Յp9p Al4�t��NQaI�F��;�/���o��bu���b���3T%z��л��m��v_��/�c�`��
�ւq�R4����H9:V�����l�vf��K���m�����Ez��)+��^n��i����:�T/e޺uU'7��X�R`�S̬�ز�ۛ�F�p9Tg���n�%��騒�o|������H�,�	Ν0��ȩ�h�q�^Q���D��; eJ��p����Y��A�|��/]�i�֑���|�����ty6��v������5���2���Pa�~�#�/�d4&K��1Zy}
V �R�l��J!�&��3�Ӻ��q�"��p�`�#I��-�˼�n��V�e>bԳ��>!���j�GD3�8��h3.��!����\~{�{�-Ϟ�1f���0"\by'�HIz��/�O4�ˌ��/*������͏�	
4��Sl�����$k�::�/](�"8�m#�=��p?����#�V�*yA����~v�UT��N�lv���5bqu�%J�07֭-zU{��7��_r���0��G��֊�����8�|&��8d�̓���tW�RmL��"}�SY>^��r��O��f��ő8��=eD�IRW�Z�s�i���g�ZSLrn���D�Z�`u@ǅ��{��h}�0�
 W�	�cX	��^	^iFiF��f�o, �"}�w���U�5������r_�/��r���5`�H��m�{5����QF>T`���7_����4�m	bT��=��"y47w��8U�˕X�b�ն�J���'�@.�8�,G@C+�V�Wҗ\�Mi�$ Wy��6W�����A8�(�{`AٗǾ�t˄n̍W�^�m���P{���5�
� ���0������	}��s'�Ttƿ<�K�����Թ��`}k2���?r��� ��u$<� Տ�c�)��[��	�,S\`P�f�]�$~��i�.����S�2��:�g{6Z�=��"�J(���&j�N�;@�ؘ��K|%ؙ�vЉ���y�Zi>�C/��F���$�I����6!���5�A\	�	�j��4h�x�_5�"
�Ҩ��v�<��8*�I�0@m���1i���*,�V!�Rp��A�vg7!c
�;��-Z|�̰_���O}���@L|�ʟ���K��ѿ%�^���vx�J\k90 ��-m-�Q�nPø�.���P���[����������n��u[V-�+�iu����F�f�n�* �`��l�|�&~ep����Q�d����5N����R��UpY��.<��|WJJ�C�0a�u�fl0�@�g&= �|���%�:�S題U ��T��h���(C�摚_��[?�4劫�[@���d�����.(dœG�!��d���Y�� �SQ-=�몞��;R)h���8*�~*����M���$�i�j��@�T��`x]D��/4j<m.�p"L���ab'�]��oJ�A�An9h��,�>.�w�Yq.*�<_��]�mۇ��h�����rp�
�Ig��E$[���)Tk�L�dcd��	
yј��*��?����5f�yP���A���Y�e&������w���%��+�cp�k2U�TI�&����0�8q-;+�E�7)W��o�O^.4�W���.�WgV85��MHȽA�o���;B�߼�]�����k��T1��il40�Xʠ�MQ�����}�[�@��[�ͅzP�q�f1Q'9����]a+��ܿ���%}��������o�����}\�@Zk�Ol�w�3��iç����&M � �4NGN����UR?���^�ks�zmz�A|oڞ��z����+A��%�ɶ�`ĸ��\��ĳDw��s7`��9=���
dwb�;#���E��������[��kM���[~�.��a�]������	Q�:L�5�lќ&g���������u/A�$Qg-{.0���*�N�^#��T2c�{ס-��x�)��<�1��.xZ�u.�9x�i
��4R��J� ;h!x{����~2�-�mMO)�nX@`�c8�n�@���!V)Ow ?voGD���)����Eb� ?��S�/b�F��X}Wʴy��ЉA�[7�� ht&Nn�`�*����#�3�J��}�u0��9�$UMcV3NN2ѫ��ި�7^]�Ƀ���� ٵcT�y����[��3�ݝ��@!e���"Y����P��Zw���rQ�hx��P����Kk���+���ڡ�`w.>䫽�?Z�n��.�N���b��|���짯a&E�SfUs��P��0�FjN�/���KU��uN�W���D����A>	����F��2�?���7�a����h%��qC�bX΀�8�1�󳑨���[R���L���\�0��*������-�Uw\�ԥN���4���H!+@�XT6�bܫ�����r1�q����JrN���W/�!��RP�P�%�ɀr�%}�aq�MQ�-�#!Ϳu"�����=��M0�B��GW1�Y[�n1������Z�}5�����2$;��h~7|ntWD8)<K@O���\�o]�/E*���ϝ+/�Ay��fSyz�WZ� �Oqę��,08T_�
s��b�jj���DY��Ő���'�>&��<��#�2%���p���ˠ�x�'<��U"��0���~�kh�КʍG'+bF��r-蓚n����]�x��=�[��fՎi�����Zړ���W��T�4���aiR)�r�����-\� 3MKw�t/�N�|nY6q<T��(ȍalڌ1��)
���}�P�9�i K�+ɛ�ǚp͢�f��A �|c�ݗՓN�x�}�WM!��!�������Ye��F��i���N���j�÷¸�< ��$}�^���ڥx�KU~�Uw�Ĥ
⒩�Ȗ���Қ[�ҋC��Ӄ�'{}j��}�
�ga[�Lv�����7��{�ZQN�)�}fi���I�$��x�:�%!"�j����ޖ�n��[*�����k�����A)hSh����(΋_��[���VsYb/k������Z���u�w���dZ��m_ D���(�ѦZ ���dQ_6~���j�������t�H�8�J:���Nz˅�����&ݧ:'T�G�Y���P��ec��97
sՆ�"�6E�hv�r�i�s���g�}��\��ɕne�ҭ|U4����I�.upcrD��~��$�<���� ӌ���L^�z�+����2�綣�7!{Q2g��E3�v�Ӗ�2+��-k��Q;J����~4��8ʝ!YɬkĲ
*�,&�=����>>�5�r�=�Z%��2S�x�}����Kg��m���\<'�êP��玥*��v�"����:�=/����=w�n���j>���(j�����!J���Qh�F�����|���A������b��W�C����D�}�	1��̔����`�bR��٦�E��K_�����믐N����X�I2�AJ�����w���n�,�₴W���D�L�> V���J���Y���=�/�!�!:�hن&�
�(WU �}��+^&���]~����)<a2���zSٗ�� ���wY(%H�:���A��s$��:���
������ߒ^b< ��È�Q�)m0~�<��5�F��
3�w<�^�6Y�jB�/������?]lv�_�]�.d<{^��B
W�ʩxÔ��{��N�C���Mk�R4��hqC�l'8����:7��by�������Gۇ.l�6b_+����j*Ok�Z�L�Y]������̖��EJ�։�� 6��Q3�O�9DG�ǽ�h����Ö!�+-
=��K4~k����]$�b�$:a�0~�]�wSa��i�B������'���!U}0���ӌ�7��7 �רèL�.븠�Z{dZY夳6��z=�}q�|���P���Q��V��������]f=�uQP���d$�_-�F�➼S���*�{)��		����LTM�����g�ݼ=� �����,����_�	,�h�Y��P��Ncd�=�SZqu�A�eS{��{�7�S��%0zæI��ꈿȢ�1�|� {λ��v��+us3O������wĴ�Y��Y��� ��.!s��=�"t�������f>�e�9Χ�%O�>`u�B�`�*ѣ�{[��v{c�2E�
g�����ڕ�(B��HT���$�5
mʏ�io��V|�xsɱ�x�97���$u��j`��������[lfT����n߂9�gD���^����K�|^T]53��w�H�A��
>-�W|��D���S%��n���pP)ѩpX�'( 7� �z�rQ̒�h�t��F��s�y������zTKP%yF����U�� �|�aL��<*p��Ro�3Y��B͆��� F&�I��;����@e�Wda�|�3\��eэ��=��o\�@5(}L�N���N���Ccs'���D����f	�%���.%+�n�S'�L;�A�����!v�,��-�=K������޴ȞO��iS�jη�50�����{�V�mŬKXOàH�9�������]vYǔ���L�`l	�f��r=&'c���5p����Z҇0���I�T�H�� B�j	���9o�ܧu��7�9�%��]��V�UH/*Jg�0�P�#��Ө	ك��e���{�;�.V�������M���\�s�{��4�{��
����7Ps��tZ5�e�~���(����o����U���3tȍ��@'w7透W�4D>����ǀ& ՜�p[�kpZg33��q	��߉��ȣCB�NjD��:�YHp^����|G�2��	���U9ߠZ�/�)��.$c�!F>�mi�CLv֙o.u�aꏺّӾ��Ds�a R�ԍ��ΛZz��8� :Vc~��W�uEQ���ſdf� ����K��>�F"V,���h����{K�}�.E�������g�c��컾�@x��t(~�y�G���z81�Z�������&q��m TK`��\����?��昢�-R?c6u���H틟)�l�!z]�sY=kA�����W���]Z:����EJ����?���c#��i(������X@&�4V����<��oAÏ?؟�J��QXo��)ޑC���!������tv�+��#���hO%;�w΀)!:j�R~<��?� ���O�}���Y	W�Lk{��!��3�RGA���=.��)�N�Bd �,Z�� c�_�uuթ�����n���F��^�i�d��C"w���Ό��Pn�{=�R��<�ǋ�n��YCw?��!R��FlZ�O#͡9����铱�X-$�4�W�u�Vހ/�PƺO��Ɛn%��`�!:��M�oXc��"<)��ެ����2�&�Ĉ�#�o���l���������&l��Sgw�m��Y��沈P19[p{n�~�}FaT c�Q0k���g�/���%f����S���̚%J6.�����f��!�x��}y8���OK~��=�	�ᗬ�F�������23�w�YM(Q��5\V���Ξ��m$C%a���Tl����T��hC�/�J�WPx�3L�ə�ľ�^4�L��Hm�ܦ1��X󤢔�ꇳ� �H0�`?�Q�L�t��1�)ɢ]�ݕ�z��#ѻf�E�_ۺ)��rD�#`��
U`��r��<�����$���~�ֶ�7�t�E��Y<(�$�ø������!����vue���~�&���4m��ur��V�5$�i"���鍋�1�x\\�u~O�����_�ޔ���M�Y�|NYe�m�V_����9�V�nไB�����yDem%D��'$=#&+*V��\�y�x����0�]�2\t���ٹ]�߶G�o'��p���/�q���pl�WG1�K#���"�[�'����ͩ@<I�A����h�l�Y��$�L��\��pUK��
�Е:p�������'�)�~�d�@vX�l��3����4C��6?��� �*zbt��a;h�ƠB/.ȋ�66�k�]�3�4�V
8Կ���;"8����hL����Vfd⁍gc�(��>��T��e��L�y%�����\�W�B �.�Pp-P�Cw�����|�ݷ�kيFq6�� �<K�q�f��f�[>ʃ	3�T߄�GK�'C��]4��<�g_�`�9�ۻq����D*s�J"��B��6�d�68�����fu�;�C���η�+�a�zc�]�h�)�q4��`f����F?X��Q��l�Tg�&(L�׏Q�&Q62G�k�C��[FZH����9>�n-o/�����S���Y�}��O�֘��M�y ��DG�I���j�ʇ'��t�X]4�骛����WǸ�9�}gr>�N��{M-Ϻ�r`���\�ù/�#�*A��ޅ�0�\O�L�ū$���;ON��a��q�A�:|�?������k�p����z�Ȥ�^wM�K"᢮kk�D��$n�~ �]	�t��NO[��J��1E�bi���P��Y�lMF����\�9&��bY5cXvG��q��+e@�P.kU�,���k�u�B�V��6�Il_d�|7��cx8�}0����^����f�tW
��m���c��8L.��lR��/�E6R��1�ڰ��k�*6�'�M�J|�~���w�e�z~�o��eD�$P���pvH�w"�xa��2l���Ck����u �X�l�N��I�:�װ�E@E?��k�����w���T� bHe:bL��e�/M!x��wgg@�x���Mf��LNE��SM|�A�����"`߳��/��SO��&D��ju�{tpP��!��œ`����6��*d�+R3�mMs;0r@��π'����H��p��]9Ө*5c[�V���N�+�x$��Q,ː���[A��^!nՈ��L(�����Mi�ˎ��%��Oe[г�d�i�ǶZv5�o���	u�Ȑ��#��<��l���#$�9&��~�Lͥ� lN�T���C�_{�2��z��ȿ	J1���Z���S�����b�{g�-��3vZ(�63�bs�#�w5١��@��
�����C�Җpz}�a�����̨q�i=D�%u���JU(�<K�tP[!�5�4p�E�Jz;�}��׋^9�^�u�"����?2`���O��þm
�ꐒ\P�o.��70���xD���4)�e{ ���Me�(���k��p�Mc�ix�Bfgya�Xx�Lۋ�.{������[+��Ԝ�Q�� ��������JT`Y�_y>�� \&�S�XQ��3q��%忙��V�Ok�5�|݉��&�1
-5�I���u����m���Q�<:a�~��u��H; ���>'�bt_�WЂ��R+߸t�V���:�=?KWR�02OK��.�
��9���~O�������҇�є�&���:�5=�<y:��4�\�����I9˚��[9"� j���i_S�<�ZF�c���諓QF�o{��"���a-Ɛ���[�N&X�k����AR�~5?ϡ�;��e����F�ox]:�o�e�l@� 2�9��i�1\ܰg���Ƿx��sWK��ä�FTH�w���� �;Kf�/^��)5�;�C���L��7ń�)�ɷ3x�����z�6\��-�&
;ej��*���p#�)4�"3�6�:w�j��Jg��#q퉼�cZ#Co�o��d8y^8�RĄ�S%��(� �8��Y�`y㷧�ww<�-�=��������-�-#�:懔^vy�.&��/B��g�@o6�
��O7�[1GB�#CFaK�n��c�����Q�<+�"7p2��o��\���P��0�SΥ&S��\��xY���m~��������
���H�Ǹk8�Jr��!t/Y}��8u���9֔���"��r��e�ޠ| ���`p�I~�B
�� 	�ђ�����r���I�3-��K��!#�{&���g?v�m��\�byQ+sǣ��}�4���Q${�I�yti'e���i �cL@�0AТ��Z���+Լ�Ӑ�� �X}��0�4�M�8�6�E).�mV��g�+��y�6?m[����?�}~'q+]�W\=Y��f�j67O�$#ek"8f��f,�`�[�]f7a弞H-z�(�I����)0�Co�|l�]�]��A�#�s�AKWe~|ߥ�x!�g
_����ّU����mjV��15
��3$"��K�o�Ģ�}��_$$ϭ�8(t����b��C�0�g��m���o�%�ŕB#��Mk��0U���^���7��J+�֑�3��'�d�s��q��
�+��lT��d|�"(�B-�:^�~����� ��� �3Q�b����F-l��ܤ W�@b������u2ٽ�Y���f(֝l& UEr�Hɞ��_�IՉ4<��ǡ1��nұ���Q�6y%����h��x��4�x��F��'K�)L$��Um�\�zd 1k��uAz���`�|'�G��`~y� 6tJϪ�GĴ>��l�����p1���"��������Gp�y�^Xַ�|�� i�Ǌt�d#�A"��m~U}�W��IU��gm�I��Ja�Y3Vg�Z��'1��j��*�o̿y�w��`���'�¸�Q�s����Q�\v�=B#�D�[G���� �7�5>�ː��9�L����	��D���{Msx* O�;wT�пO-�4���'��dw���-�����$��j��<א{�B�wn�^(^�܈_`i����s9�`e$�c�H��"lu�r
&>�=lN�0W7 c�A�����hv縀�`�8����]�XU�D�>K�'T��yeO�S�<�蛛������� ���:�6#�q��诇��1��}��R����9��Ah�<��W� #�U��sK8E��ߥF�!x��	�q�V}����/�z�i��,0��q	!v��:)v�����^Ƅ�x\['+Ɉ�8ꁀ��9�^N9C�ń{�ҽ���8�q&V��ńp2N��|F͑�̷j�C�(Ȧ/�Mu���x][{��X���S�pȮr�(�.2���:�W�n!���8���a;Ҋ�wMڥ��->�'S��4�ϡ���}�H�dٻ5�MZ@�Dd�}W�"C5j�*w��	ʮ8I���@Oθ���I=�T�He���"���V�b�i}Y��4?��(L�0\�^������a�;�{(&�\� �ï��+�� ���hX�f�.���r�m�:.���ҟ2��{r���>-� 
"*���gEoU�~�Q6�RL3��W�P3 ��}��n�Y��) v`�k�9�"~S���Ÿ��Nt.�� +��1�n��F"���e^�%I7/>����� ��z&
L��˃�D����vXnF(t�{��+d� ���74�������Q}\�"��%3|G��� ��7t��'ڭ�߅q��Q@~�����g�?�c�kE��˒�-g-���V5Щ����J��H3�U*�ߠ۱�c�ֳ>�^k�" P�MNz�5�3���e<�#�~��h� �������wfVf�� ˛�_����>R��d�1���C������m2n��� �挗+����h'kA�#�r&N2v��vDq�"�-Ӏ�&�)���;!��������~J4�|�GxipL�������6v[�,-�rN��.=������%����QЊL����7/�RI1�6@��H���@�/��
f
���s(Q�����T=m �=��\�H��|�ȥ���� �uq�00��K8��SC�͏�} ��L"�wT��Sy�R�09[1�4�5�ٮ껦�M��Q8���
���h5M�!(�-t�iH��L$�ʊ��C�
u���T{<i��X����y� �wy���rn���A�-O���ԟx}hu��oa��iUWLe�=+`���Ⱥ�~��oC�bH_�<�?�i��$�1��K�L��5�m�rف΃�t�*����E#��Őx�{-|uT�Nw��c�.7�4�|Kߠ*�a3���*���1t�M������u�
����p���r^�0�D�����z���7#�s۽�R���+�ߩ���Ґw���%��،U(!�Y�w�V{�����=�Z�L�d ���v���j}���Y�4^�'�s7��=wHZmvamC��e��K��DJ�36�B2E��e���E���3���%[�	�c�s� ��n�Y�&F����!
b�]��S܋���/i@�~	hsv�{�!W[늩.����S�2l��ʳ���Y��Ң��{{��Bi%��d�e=���RE�Д��	o��źԏއ�t�1�翄�Z�^����_��^'@@�-/��Ϯ�ɏOb41�!����ld�LD०-p�OB&r[1�M�,3l/l�_��Y�^�)a��L/陙�m_X��,�S�;�Z�=(	:~����_ 5��^��B�|��<;vz�"<t1�Ȳ[����ii�lo���<~�s ��4i}~x���%��'�?Ɋ�����~T�R���K�0�y�`������V#�h|��S�,����!����%'2�U'yOw�~��4b�e���h�o-f��N�xH`���� �">�9L�<��K4f=�;����4T����R>��r���j�a3��.�����(F3�����^ǵ9t�Wy�+��zB4%�3����D�����K�:_;�2GZ�b�^r3o��%,3��~��lb���=8��L����3��J@��B9a�������ܭ>[Y#wOo�-��(����l����$f�y-�>ꩼ�s��v�6ԈK��rP�|}5�ײ��{�������Ӿ/"��Vj�{U�+��>F~��b�h��D}�,�+��>�,���k�s[c%$�C��}(\"�<&��M!7S5zT��!Z� pwEX[�S@t'N���	�-Z�W�"H*Y�cp7m�ߧ�bA�-�	A��{�x�s}�҃m�NE��L�4;<c�j�(Y����|���QP-�Uy�H3qp�j��OBu`�Nw1�II��=,t�����������/;E�I�	���Ђ��ڙ�Lٺ�����*�+��qۦ�jg���| ����`���s�ȏ���B~���͕�x�'���ׇ@c�{���w��o7�7��^�I.?*(g(�z����5�HB������0�,7�q-�C�
>�7�h�ԚU��cA#s�`'�N<��J	��[��~�*dݓ�m��r@夼��,�|r\�H�7�0�B�,��ܽ���iT|<�
��y�� 7D}���09m����2ח�n}F��3rs�$Yf��C��(9�3ך�2+�&J`喃7�n.w�7�j��&���R�/�[���L��SG�x��_���>cgrd�4K���}P���%����0�E�D"|��H���la'�kؿ�U�<[�j2�шA0����|�����΃����ʉ���)�<!�ӮCd&�9�Ӷ����1_�<�I%�ZӖh,a7�XXawP'��seӮ��
��M�l�ǎ(p���U3c�֔c5��C�0�v�������rIW�~�5� ����6t}�73�M�QOv��������l�׭xH����_���Jl�䥦8*�j��;��A�j��s#t0o�{Ƚ���G�������)'��4i��lR��/���C}r�}!�*0���*�c�вf
���J�ST�)�^.�gH7x���s�K�.UL%�E��8HNp�Y:Z.9��	���hB*TV���8<
<��8�xY���tT}^����V�u�FS�{{LM[���S��͈��"*�F�($�8;uw��t�R#����������s��b���]��T��
ff�z ����k�=13M��R��:��c(6���-�ٔYd5c�yi��doLgVeF��HƓYP�Id��dJ=':�����p��6H�:�lJ��-�e!\A#YIA����wX95���a,�uA! `���q,#;%�*uL'���-� ��҉�t����Cx�u�r�m�<�C��^���o����6��AҎ��ʊ�Y˪��t{���k"�7)�Xwx����'�S���1��C�m��vPҞM!d�:6�qu#��q���0���	&���0��=Q��_�w��] �CT�y�*u�՘�!yt�$�Ǐ]w�)�,c��D��U)���c��/��.�X�Q6g6��׷	�d�1hf[K���.��΀�MA�x�p^JE�Z���8G�#��!���1�;�:`E��ؓ���z�Q�1��VX@"�����ʐΰ�b���)�)��	�	R�HǼM	j�)��xu�H]�7�&�x~渍;y ��'����L�UT�������A�:+�:+��a��Ņ�����;p%���p����[=�+m����R�D&�� ׈����s�9�uȇ�@�AO�����\�J�=�-lq�`A��X�>����v��wy��~��e�FH1��1�w���y�lA�7S�&_�y�K��dN�G�("�~�ę�u�()��V��]��³��I���7,���ۊ����S�cO�G��������[�\�z�XG��7������P�a�]��H�i�f��B��N���[̸��0j����O	�PNz���	���2i��2�����gMX+����?���ό�zL�0{U��9�1�C9�ɞd/xJCi�"�0���cӻ�:���\�L��������bW�^4���B���:���O|J���Nm�9o���e��jJd/
3�`��-{��FQ;޹��&�v���;n��4q��L���������;S1l$��w��My�٘�'F��Xh@��xp|�/؎��4�/�S�����?���+c�#����U<o^���e�8�7
԰lyn]�-`�a�r�u&�mY��~�L�wo���\�����sӃO���ã7��`�8��z���Lh��^��o�[<��٠��!��e��}��>t? ��(��coW��_�O�4�.�EQ.�s#�/XT���4K�j@���Y�������CHC�e{��&�R������1�xX��"�x�^9=�+T5��rw��l�^�4�tbG7s��4W��4Lt�м��ꉮ���0��>�,��5jc�i��!�=��������ݿf�ܨ�Wߺ��.�LbBl3^&"+��	�f�EH�lTt��_�S=�S��!]]$q��#F�}�%�`B������<������L��Ǻ:/��]��e��.�4-�3�?�+�\Ņ���a�0|^���Ŕ��:��_��L�ئ�,N��-�t+_����{8*, e4�d��,�߇����2�t>�M�tc��=����!9� �����EO��-_O��O�ߟ�_p/f8�����2�x�N��^�､���&�.4ѳ��	���?<��B�֪��:j��U~ڏ�&���=�їE*Z���L��di�P��5��W[w�g'<�!\	[$��^ j��&E�H)�#������=�����V��rY�=�h~�6����pB�DИ
���#>;���dhvh���r�Aj�a��>���5��\D�nX���A��B����xH��B������W].|�j��+��a��Lv���M��%��Z�Bp����s�q���!!8�g��
�X���B%4ʣg���~�]婍�g�7*(��-�&��G��]ozێ��՞>!3-�᳡hSd����it��	��+;��in!��:�0�H�r��=g=���/���0��1��mR ?�^��z^$�69�P���1�D�
!W�yqBMx'�K�$��}������%�RtZ;lM6��Ћ7 �4Sm��~�.^��J5+���ߏ7����������)���!�U��PˎjQ�m٣N�@P[�؝$;V��d��NkZ]���!�<%C�;%��w>Uz��~%���snCT�?�a�#��W�Q��^��td;��1�ېG�*KKz_?G� ��b"NG��&mrlZ\G�\L��Ɛ�6%���4�2��h���M�W�R� �� *�n;�]}s_�����/������7 �(1��sS	������֙�����u�t�tkWbߥ&2��ry%DQ�T`N����+��r��_E��>IM��j�ι�_F�Ƨ\=�M"���W"\�0���'�o<�pOmK�������>��Fs������3�hv���:I����$E�{N������H/�?+ ���(Ly�E���b�}f�z���x�\��X?���@HzY���dvLrD����"T7����Y�Ą܏�!�~޳W6+����M.��q��<����%c�`��q����_6��y��U�,3�xU5"�� ?hjO����zPR���2ǽ,_]������<�,��JW<��1��R��+���d��( lm�p���V!�t�ɦஂ����KGO�?�Ux(���\��X�d��_�v�]5_�fM̙)Q�r}=�)�73���~d=j�c^R}�rX]&�&���pk@S Nz(�G^9��G\H
yF��:�"v�� ��?�\!��|;!xc#���k��6�X�	=��o�Beܕn���_���c�j��tIB��[ܵ+LL��~Y� �F$�����ب �YT0�<Ae�Q��l����_>�R�E��"��0��&�0�u�ِH��+Ӊ�ObJB"��bq�h&О��%�(\������m��<L�k�}z[(��O"ў��?���1?iw��[Õ����C��h��(��r��=AJ`�՝����#8NJ�g9ف����%������Z����B19 gO������	�7���xh�X�k]w!Ӕ+�;Z)�U��;�τ\��zei{@��
��m��j4Bjl���S2;�垟�����9&���
ߡe]C6�f9�A�$�x�'CBǕ�M����M�}uD���&,�we�$�:q�iM���n�d���Ϛ_�O干�D�=l��nF5��~,f�e�v��WE�Cٚ�?MA��N��TҸ��k��ot���a�4>
��B�+��Z��XO�<H���O���^�>��'����,�Iy2F���=ߘD��H* 8�d�����J�(wl���${�n!���xgt�����7)]Us�،֭�>�dl�kb��1Z���9��z�.���+����{?y���gbJrbx>3����?G�DM\��]^�q�t�g�?R_1b$�J08��#)u�N�&Sw#�emX?����<���$3*#�����V$�<�@�m�N��M����Y�2}����-V��6r(`ڱ�v���$	����1�O��
��{�j�=Ih���b���q��a&J7�Ǡrگ�<��Mx��-�>H����ixHi>J1�[���t��AE��Y镞.�.QM?�<n�y��.���ı��*c�J��g��$�<Wj7:G�F#UJ��bS�[4��L����D;ԭU�*�:{4k)b�K��"����.9 �9��a5�����;��d����z'�9�>���Z�:�DęB��XŠ�\h
w.&`7��8��||��:b:�����3�<ڀP���2�>�q��KvҨ(��}8�N�����4��s/�k/dA��GU�=���ޮ����#)t�{��r��R�����9=����;��zd3�"��k���O��@����k/60twok!��gIb%��bݜ$��a�O���:���2�6�U<3Gɇ^�χ1#^l)n�D쒔c�j��vto����_��-�Dg�^��OE��]������pkz�2w`p�	תZ�u��P���G�W��-D�H��A���ځ�
G��g�c|%z�XBY���toڼ�y���u[aC���{
D��>8�'�1b=`��T�q�>�3�+�����T��>�#�3ڝ������j�s�i��"��=F�!��3:��~n8�ֻ�EF�'˥��{<���0^m�}�	��
���ksQ�J)7�J_�P۬��-�7�}�΅0�ٲ�t� 1�t����d^ ��b8��翋��q�PI�@���o�}��%J�&�\Z�\�"����Ji�����&o��2�QA�դ����1gd������@��f��;����ex�=*I��^����nOÊ[���G����'��,�G�����"���ou�+͖)~o�SȮK��~V	n�s#Q��|�����h�r�ʮ�b�ᷱc���htI4�H�{@i���ѵI��w{�z�o�Rg\V����]я�S�o=��d�:56���]33q�#:g0�vH�vՏ����D��n��9��F�p��Op0X������M�Y�v�Mx�]p���jaLR2U�w[S�"=;����iV���}Q�j+4J?Q��7)�	;I8PF�B�V�Ob�gu8�*��?-�����eF���J"3�D�88�55!��!, qe��8%ZvY��;�l�Yzhpm��1B8Wi�U�ܳ�O�H+���g[]�[����.h����g�8I�$��8{�e�x&��>@��n���+�����.љ�V4�Gݧ/k�]���%e��E�����H��n"�rI|-�8G���-U]���"N����w}�;��}�%�!�K��;��""(�9��ZИ����m]f�%��a磡�'s����ј'��"��0���4��K�[��]��M0g
�n���:���[�6�Y:$��Ǎ�uj�P'L1�B��$��U�tb��nSQ6uQ_Т�Y����?VH�c��4Y��Iu��2XuY.�~b����&B�Z�G�[��h94/!nқ�1Rq�0��� ���6Τ�T��縖����52��u��<�Ϥ'�ݔ��:Fg:#ft�WVFm8����n�H�d&����6=�	b%�o&= �r��h�0?m�㻙!��ӹ�"s�G���T&<B�7�qt�g�����2��l β��:��1�h�|�'�h;��`G,��K3kh`�c�q��L?��y��SS���'�O���!*]�a��!p-[��+�qM���&���������I*��Ü4�VB�'�'�10k�ɟ�B���28&�$$���|J��e�L&T"�7���Pv�uko�����:)!q-�[YTB�J.�:}RՖ1��y]���p	TZ� ���,�	TK�Q-�X�c䬫b�⻠�d/op�5�C� Jx褘i2�Y��a���~�貲�4�t4	`Wb��RI�"�vU֫G�΢�2�����gu�b�%1�q�_��t�^Jx��Jv��_6u#Jv�=�L;�d:�ڳx�����;��E%�BG���$6�QGr��mW�=H7���2%"�.���V�Z�+h��LI9ÀZ�j�����4�˖}�\�&6��&j��%�s�Gٍ��Q��x���ڔ� s@'.�բr��s�76��[炜�/+ ����=� ��ණ;H[�z?g�J�i��r< Ȗҙl�T�b�J�5͇��KW�w����3ԍX�%A�ӡ�N���F���fD��Pi��ξ��r���a+��T���β�\`L ����E�UI��O�����:P���{�շR��	ړ�1J��Ĭ����c+� W����n������!J��p��Qdع4g8d�B#�DzI��~���ڝ��>�26�>T���[�f� q�H&rz�5�/q�N���Ԟ]@_��J��Rw�r>n��|��`�2#<l7N�B`1�#�a�W|s`�����ZVr%h�^K��⤲�殶��7yθM�/�KǏ�ܥ�{k�U�)�V���"�$�6[\�]�I��e�QPޝӨ�˙|�K��+en�S�E��,�f8K85�e�!'@M"�j�.�>zʳ�Tr�	���޻�h�M>���=�����O����r~rn�N�Z,��d���#�xHp�|�`�����Z����K�2�,���CH��*��'�!�]��K{&�j�y��Q����(��Z�Z�^9�:J�R%[Zu���-�椊!�3DP/���V<N�P���Ɣ�����u$s`�������5Te|ǧķ4Nev�Zr�����������LUC�rth�z����WC	�ҟ��2e@�c)޻Śh�Q�3ӕ�S��N��m�-S���E�� (�JZ5(�� Ԩe��)���u�&Љ�sʀ�(�ly={㘠͖5�V�=�Ԍ�,[-��e�[C���.| �AUu�	rEC���F��Uf���a�%����S�Z�h�5k�w:��]mfkI��r�`H�ɉ����J8R"��G���N�h����=J���y}�U�8e�u��[��7��׍���c˥�Y����:N��H{�";cw,>峱��m�J�. ���c[ܭ�ß��u�\%R������!W� �EA�Ȼm�%�����_&"�m����[T����K���Eyd6��@��S�N�o�n%�vγ�F^1�`h�!>�L4��uY�LPS	@T�ϥ��u\D�Q���)~@������ڋ k���3��\�f���ŶH��l��sk��[4��|�I�u��� �ܩ%!k���vf2�(���I�m���A�&G��Ӣ�B=�%��x�'�^G��:霒uA%u��}�
"���M���}IP��Mi ��k�?����^����J�!	��4�ajc��j���lO��%؅O�:�[-ZÂh�&�BV�_��l����ӠE�߿�z����*{��1w�$�yj3Ϟ��ܖR:=�Vӝ��m�"���}��d�N��j7�f�;ќ���c�}Jz���P�K�b��R�=�!@��~����(@�W��Q��[(:^�jժ�ĀD+��шfމ��a�� ��fuFJtyЀ%��%�A��h
��(�U)tA7�)Ħ0�-'[wO�T��f�H���ջ�mR�S�i/��G<�
1�u)c���u`um0z	+�xa�fE�3(�B�}��AO�/V>ܔ�Du�*ny��ȑ�(S8ř)��.�&H������RN���!5\���� ����>'������Տ��g�R�/��7��-* "F�N��ִ��{�7��.�7�"17Vi���A8z�ޚ��	�����p�N`K$�m��Tk0h��e�Ӆ�ir\�4^�5�/1�?1�\�t.Q���BQ2�^3�I��*Jx�����<�!F$\�S��_>�P�	�A���/�f��,������2�fI���a�!0v�Ӧ�((��}��;9����f�+�^�58��Vm�@�Vf0�i���/��Hm�|�;�]�*G�v����aM7�y�l�IcS>��?F'��dS2}���h��ຨ*�goV_��p�^|2P��kp��ɷ�hakJSWr#��0�4�y-GیB�S�'7�����1^�pA9=f1��9s�u]�|����D�XG挍s��ޥ�xj-�*�+xM�P�����5<�Ma�w�	��n2�ҷ��������e?�Y]�e���;��%�Ϊ�Ê�JD�B�'͗����@l�{X�\ �"�}a�����ܼ59%� ��9��x�G@%<[�Q���\����ŧ�	aRX����Po����������V��K�j��SC��V7��(x��bpl���y�F�3Sh�e���Q���y�R\�z���z�i��z8��Eׇ�U��$��x�Xu��^K���=�M/N���1�b�p��V��P�P�U�(#�jV2�5��^�u���M$OL!SA3���yto�מ ��^��P����꫗H��x��b��ϴP+H��+�w&ꐶ^��=�c�aH��$8� �15zQ��tR^������8Pil	y[�ϣ"]�����q!��,M�	j�g�����sĻ�<��<[��-�PƂ��J����
��9?=�z�pi[%�NQf��������ct��q�*d��U�S�$G�;�oD�M/=�$傘�<TX�ŢD���<=V��m��.���qbe�qϸ��3�\�&V!�y�?ssF���f���H*:%+�]:Y`7-݉뾄}�{:-*8��qIw�ʘ�:7'�qQ8�ϴ8��u�� �yWya�/��ͦ�^n�&�T�T�#���mh

P[dҘm5�.z#���<6@3ej��@uEP��J�c�pB�Pu
ٟ�bJ(>J��C\Yb@���信��3��Ѡщ����[����(ۈ��j��N�J5%ii��~%�u�����@,>W�K	��Yڂ!�^\YΔO���sj���^�i� ȃ����2��O�/u���-Afd�i�7�򛡖H�L�$����a�6��
xٞ��x���"� i�=z����o��=%}� J�w�![~�>e52v�~w�#��ux�Zژ��؛	��4�EjL�	�T���J�>�?%�_�L�Oh�T��8��6���i������7Ɠ��<�iI͉h��1�i�×����3A���=9���
?c`İ?�TZr(�y_Mg��Ɖ&>RC��>��!.�44E���젍��Cc+.$g���y�HҾ�V�I@c�[o�<�4V7�9Z$��6��+��;����9��⿯$��t�y6�2�!䌙��_Tj1m	�U�{�����R���ѝ��a�x��V�8�����6�'5��7�k@�N�D�kuKAu���@�A�yi�4���OL��D��'�H��X��8x�G�{��:�7^��� ��*h��������w��@.��Hc}2p[e[�o�ӕ��礼�3��ï��R1�s�cI���&��q��HU��˙���RE11� �c��w���	HK�xh~C1u-ajMՒ+�imη�?@µ!�I2�d���Z���ȗ�>O��G��v��`O�5 �&��Ȃ�M�S�������;��]���')ϭ?�ia:�
P��"�'b1~�M�;`N��_�gbl�%����!�P8�f����Ӆ�Ԟ�E���%�Gu�Pێn<?b@��~��Y�F�?mhw��)�"�hR,@�LxJ��̇����=����E�����d�xp�� L=��K�?�M�q���4�l.9���B��H��>����{U[�Y�gt|y'�J��h��iG��hl|uu���E��M�È�y��^dN>��S��Le�mB���7`g�������]}�\�Ӎ�	Ѻ�%�,��XB��o��(������լZ���u�HL��a>��L�z�ھj���z_�`"3U�	�/��#��S�"�Uֹz8���ᐝ^�J����xe�՛���]�̧�BG)��n'j�D��_�ҞP�$�}m?�uS�q�����-��0t=���-��Y.�_|y"4
��8�� �;��[��xn`�a�:w4���`hy��0�%�g� y�DK�p�Z�Z�ń�4��X�I�����!|�J���E�D�b��y�lZ����c.��,�KGxs����?�b�A�v����.�HT�r_��	��x���ͼ0y��&ݺ��Jۍ�<�<�L��`��5�q<L��6�!�_F�ԏ�J���~��ɷ��Nr�gK��`h����hL�W���<�����j	`)P��]�1��^�6�� ��p�J��۸'�CM��qiI ���5h��5������J/�=��RQ��/䠁h �����C:������CŌ�պ[�g��t$���-5Y�����y��Q� ���<,��K�P�X_B��_��?1��DZ����"����ϞŰc��P\�h/9g�$��w����x���A嘎�1��mUW�'jK�tJ٥�����|�4M�5���Wfb�'�kDʉ;�{��FE����J8��Q�]D����E��^�֒��l9	 d?����ո���*�`#�*�ǜ.0Ս���.{w l�E5�Oj�MM���A���?�KRXg^kU;�lO�_�`�eЦ�$ZTNk�_2e�@�ܼgp��>��?.S��"�GǶ!"�Z�cu`:Hl�kd�dU�_�8�����%3��$l�h��ܸ�n]�~��������no��Lf�"+R��U3��`�W�I���؋py}+#�<�H�V�y3׮�y�@���04HU ���k^�T��7���6+H71>���>m��I�O�iy�����v��9r@Yg��R�׻���p\�G�ya�sE�i4���*&V�Oy������m�1�0�r��y`�t�eY�P<iI�n5\K�xj]�@���?��D��v�zc�~����1%�3�����Y�C;���L����́Q�ýJ�[3�$���9xE��9����b$OV߮|���C.hDI�j�ns:�B 2�kZ{Hy��n�D#I�|�[$�|�&�1�ݢV��OO��.3���
��DC�^���!Ke�A�!ԩ�xM*P���]����`\FVrH�x�j�U���� p��)�.�!lEt��cq�,��]盐@�e���~����bRmˏ^]������K�b�l?�Ѐ�1�������5x�-�����!|������o&���e6�a��T�u����K��{_o#1�_�;�a��4����=۩(��\NZ�/ܟw���²ܡI�@{cC!k�)��NLss絫x\��a8��}k�D#+�&p2��\�����J�J(<i����vAp�$�W,p����A�",���{Ɩyq6y	�'�do��n*���&=�K��q@���/"�~��|�l'���=+������3�!��� of
�*����ƶ�0�b��+���/m�iG�n`a>K*VK
�2`5�����e��#�+��lAʆ9 �n�1&���Q䝌���
-$�%iaZ(�u������K�Sa{̩�m�Q���������kִ��t���E����2([�JG[���1!���������:N�@��z�*��L9k*w����:7��ֽ���h����,��)4gl���zʎ�Z��Sὣ2G.�[qN�l��*���?=����]�����>ݾ���C�z�<V���vȯ"�$�/�4���4�vI�`�4���VW���`�qk�HV)IL�%�X��l=�T�_'��lQE��ý�]E��a�I�5	���e�=e�w�hNնJ�t�z�4��W�B3>X;��f��Uة�(���w������Q��	�3�+'�ò�\�I��7m{�#W]�XN	�ӎ��k��P�wf3�C��c�W�A�8��;�R�K?�_G�`y:(�n�<�KƔ�fBr��w���O��@�;`�s���OXV,���� �� $�U�h��M�aE��q�7Z�m�w?�WK�Ӂo@U�M_`�s�Q
Y'K���U��,_l�I�h�G��L�E-��!����A�U����f!!}�D�t>�-A���NP��_b\������7�x2����h1����?D�̩s���&,�E�4\ߕ��	�J$8	�]jfR��;XÓV��{��`�bmRF��@l��R�5�*�M*o�0��ʁ��G�K�&^����]�5u憎�6��y��w���^N���}��0C�����7}N������/_F�;l�ڪ�ѕ��Q4�T%K������%��騹MF��0���0koo����;1>����\
�7(
�q#i�Orb���.nWl(���!�g�n ��PK�p�7w���o�<:�{ "ث��CD[H;��C� ����slP,H�:8]m���cdԥ�q����2�P�V�'C'����4�f�W��'� �Y3���F��LԯU����z�Tæ%f��5�%��ԭ�
6�`�um'��0�v��>���p����� ��q	��6�[�41�e�V��_v��T+�]�ef��ʡcT�"�-^��4tn��Z����h�e.�}���Uqmh��G��mk�ٞ�3}���m���{��*t�«�2`"m�����^�V|�m$�����,��gt�&o��Hޟ�"�h}�%��+0�K�}Mb��@�RsBt󗍗��̸�5�E�U�~1"��fzn��&q�ݰ(�>�3 ��3�ռ[~��F�}��=-��:�v1�ཨ��\�(�����>�����E�
�^ӥN9��cH�l�a����
<\��e�|E&b��0� �cv!0<d��$��!6�"� �<@,�	L(C� ��*.�}�� ���`s�;�w�mp���(A�X)huM�?kD�d"&md+Hѝ/�����8(�y�Ԯ�Js�%,�Ͳ��gK��9>�B�����w/#ݸf^�DU,���,��"*�vJ
!<�f��[�x��⻚�7�x$?�"^��^ǂ���;�UL��\�]��S��n(k���};̥�h!�9Z9c��iHU� �%�=CeNYG	˶�X��a(����{!�k4�r���	�oȭw����Z���
��TjH���u�N�O��ƻe*׳��A,�U�ۄ��.c�ݰ�s?�z�]E��eg�2{Ċ�!�<?|�Zz��uxa�8�}E��`'.���q��5���#R}���Ըj$��W�X,U
ԕ��(8T��ܑ?|��?��~��wi�����c�'S\F���j�_s%� +Ԁ�6�q\�4e��鳀��z�O�Е"�NeY+��í��$�%	�5H!�����96���@�/4%���'�'i�[yJ�$/G\�4z3��+啀��������\��2��T86�j�t$�B,�2����	O�J����|�ľ*���>a��Q��O�T�������/7��tߦig��l�[���K3}J,��e晴���OQ���)ܤƆ��v/j�ֿ�Q�=PhK�01f����o�6fL�Ӳ*�>�V����0 Z.xwn0��֞miD�h|�JbC���� �aQ^G�Y�� ��|��a�S���4���$-jT�F	�$�z� �/>�����%T�b�~Hrk�%��*$#~����_��x\A�
"�K���wW��f�8����d�A11̚i�]]N���p�,��ݗ��CO��0��~�Ep�*��Wǩ�L*�(a9K��*�X��'�$�������؊��|��H����'�;o�gnV��Q���{�yB�� 6��0=��%*�����C�<�د,B٥Ι���@.�CU��'�3y«[،R�S���[W�Eӊճ�e� ۼ�h�$=w2�P?2şԠA�չHm#��~h��e��Zq�|.ݟ�;����)~Q�@��HX��h~�=0�=s�����aZՉwL2/�L�K;�apl�����������K��l��7�X;���s�6�W�5}�|צ���ƒw%`3G��r��^��:E�"��b���C�[ ��H�à��G�k�����������Nڽ����҆e�b�� m�"�c�-5b�W1��z�ݍ"9�4\���p�,i�b�,�����'�m��1�#����۴!6Gݮ�._��A���v�I�%k�P�zx杘��SKX�}��_6f�˲{�����:�,�[�KSae_b�z������L�-���X��J܌��a��"�ɹ��r/�Ю�\xl��X.��0�|c����Ť����*�>�[cL�Uv8���El���D���(pҞ�_�~��:j�OaO��2��9�$���X������z-�1�kB#t�]wn���dEX����΋T�e�=G��T��:�r�&�^�$��\:A9'V��Gz`b<z���J��_��b�� �{>BH<s���;��ɸ�8P9 7*D�ޑ�{�*��*�6Of*.��]{��� ����e�*�k�����ť�v6�S��4����'�;8��Y�}���y��CR5�Ћ�i�(�)���ƺ��qP2t2ɸ�������|էX�2�����E�*ֵ�
ۖ�MXI,83�`������Z3���QX��s:�s}f!$N��O:�V@�h�[�n�0��;\,I�]���c}f�hD��[w�;��I�m��Y�͂�IH(3���{�k@�`���b�q���0�u�Ό6jV:��d�$ Zʒ"4$8B�rZ��:-�:����m�+>��ږ뜉�ݦ?0{����kԨ�i����F��6Ac��qXD��=؇�v�-�*����y��J(�e+��i����Ly��(Z��L̀�~����{v�3�)+_�[q |R��%_DjG�k��qIg�y�!�_�G�
7���3''�cC�(i��A �?"��4���T�����{�m7��4-&	]�����u��C��W�[��0�.� �� �PVA�)�3Z���O�A
_�q	��9���*��uv�c�rF��q�����z����^�H�8\\�`_dI/�6�5�sc�*�*�ښݾ����@FF�s�D�"#:���F�ٵpl^��x��c���8��D**���3��'a�;'ʣ+7i��YMS[��0mB'+����R���K��,�<�36g�Q#>V�O�8 ;h��h�2���k`�]�EJ*oY��o�Qy'�ɀ�!GQZp���˭H
-G#�؍uAd�*�E.(v�Y(t��qLɖJ�b��\��"Aeڪ�g��YzRF��>5	���"�K�,\���e<���9g��`�#=�u�$��_8͘S���3�x�"Gm��
p����/�Oi�}[KN���Z�r0�B5��S��#S�HS#�ˇ�"qE)��"���(��"�Ae�S[�a�ٙ1O��6���7����ش��+����=}�
o£r�$��#h�Yd���h��ĩ��AEC�|�e&okw&{�2�WM�?g6U���U]ETw�Zf����]���PW�6�% z�,'ksʵ,D�,�Ç:���L�q*݇*��_�����71�z��pp:���6�=ǘc��kc���3�O��~)�ӾH0�wx�\��_�9�XV���W��׷����TG*��P�\xX/�ّ����ߖ�U��n���BR�A�dv�=.�]����5�8�_�m{�=Z��ws[����XY�1��.|><9�~%��d�6��pJ��۱�+k�����'��流�v��@����T1��� Q��ڡ��&#e�)�ם���6�ɉ&�֜#���tʌ�}�4�$�:���4b�P�-X!�ϯ[�xb�Wm Sy�o���4ZON|��"3�)GZ��!zq>�2Z �=��ާ)F�.��\`4O9��O0��ĕ|����ef覹�7i]�݃��c�X4�B�D���i��"e�jТ,A���T}��|@�3,�AI��p�8�>	:�����v�P���}L��8E��0�09M�ŦѦF�s'9϶��-�y�go�qu�F�
W|o.�x0�U��2�5��sf%N��䐪>��3�9���@���1���7��(>F�����ZƬ�YIL�x�+=�79f�<Q�Ι�8N^�&`O>N���u������T
�LX����a��&�\�6Q�e�Μ�	ep��҅��M��< �)x �N��