`include "Channel.svh"

module OKCoreTestHarness (
	input  wire [4:0]   okUH,
	output wire [2:0]   okHU,
	inout  wire [31:0]  okUHU,
	inout  wire         okAA,
  input clk)

parameter NPCinout = 32;
parameter NPCcode = 8;
parameter logic [NPCcode-1:0] NOPcode = 64; // upstream nop code
parameter PCtoBDcode = {NPCcode{1'b1}}; // downstream traffic with this code goes to the BDInput
parameter BDtoPCcode = {NPCcode{1'b1}}; // upstream traffic with this code came from BD

// soft reset, generated by okWireIn
logic reset;

Channel #(NPCinout) PC_in();
Channel #(NPCinout) PC_out();

OKIfc #(NPCcode, NOPcode) ok_ifc(okUH, okHU, okUHU, okAA, clk);
CoreTestHarness #(NPCcode, PCtoBDcode, BDtoPCcode) core_harness(PC_in, PC_out, clk, reset);

endmodule
